** sch_path: /foss/designs/ttsky25_two_stage_opamp/xschem/post-layout/lvs/src/two_stage_op_amp_lvs.sch
.subckt two_stage_op_amp_xschem VSS VDD IBIAS VOUT EN VN VP
*.PININFO VSS:B VDD:B IBIAS:B VOUT:O EN:B VN:B VP:B
XC2 net1 VOUT sky130_fd_pr__cap_mim_m3_1 W=25.5 L=25.5 m=1
XM5 net2 net2 net2 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM6 IBIAS EN net2 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM8 IBIAS IBIAS IBIAS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM9 Vz Vz Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM10 Vz EN net3 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM11 net3 net3 net3 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM13 VOUT EN net4 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM14 VOUT VOUT VOUT VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM15 net4 net4 net4 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM16 net2 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM17 net2 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM18 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM19 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM20 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM21 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM22 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM23 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM24 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM25 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM26 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM27 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM28 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM29 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM30 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM31 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM32 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM33 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM34 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM35 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM36 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM37 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM38 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM39 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM40 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM41 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM42 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM43 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM44 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM45 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM46 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM47 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM48 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM49 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM50 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM51 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM52 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM53 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM54 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM55 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM56 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM57 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM58 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM59 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM60 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM61 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM62 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM63 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=3 nf=1 m=1
XM68 Vpo Vpo VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM69 Vpo Vpo VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM70 Vpo Vpo VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM71 Vpo Vpo VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM72 Vout1 Vpo VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM73 Vout1 Vpo VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM74 Vout1 Vpo VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM75 Vout1 Vpo VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM76 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM78 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM79 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM80 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM81 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM82 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM83 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM84 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM87 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM88 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM91 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM92 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM97 VOUT VOUT VOUT VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM98 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM99 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM100 VOUT VOUT VOUT VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM3 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM4 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM7 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM12 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM64 VOUT VOUT VOUT VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM65 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM66 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM67 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM77 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM85 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM86 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM89 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM90 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM93 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM94 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM95 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM96 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM101 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM102 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM103 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM104 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM105 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM106 VOUT VOUT VOUT VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM107 VOUT Vout1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.4 W=1 nf=1 m=1
XM1 Vpo VN Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM2 Vout1 VP Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM108 Vout1 VP Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM109 Vpo VN Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM110 Vpo VN Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM111 Vout1 VP Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM112 Vout1 VP Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM113 Vpo VN Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM114 Vout1 VP Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM115 Vpo VN Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM116 Vpo VN Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM117 Vout1 VP Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM118 Vout1 VP Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM119 Vpo VN Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM120 Vpo VN Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM121 Vout1 VP Vz VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM122 Vpo Vpo Vpo VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM123 Vpo Vpo Vpo VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM124 Vout1 Vout1 Vout1 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM125 Vout1 Vout1 Vout1 VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM126 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM127 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM128 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM129 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM130 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM131 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM132 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM133 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM134 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM135 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM136 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM137 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM138 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM139 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM140 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM141 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM142 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM143 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM144 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XM145 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt L=1 W=7 nf=1 m=1
XR1 net1 Vout1 VSS sky130_fd_pr__res_xhigh_po_1p41 L=14 mult=1 m=1
.ends
