* NGSPICE file created from two_stage_op_amp.ext - technology: sky130A

.subckt two_stage_op_amp EN VSS IBIAS VOUT VN VP VDD
X0 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1 VDD a_6939_14134# a_6939_14134# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X2 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=88.74 ps=647.96002 w=7 l=1
X3 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X4 VDD a_6092_17969# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X5 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X7 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X8 a_6681_4767# a_6681_4767# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=18.56 ps=137.28 w=7 l=1
X9 VOUT VOUT VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=4.06 ps=36.12 w=1 l=0.4
X10 a_6105_7756# a_9061_14046# a_6939_14134# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X11 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X12 VOUT a_6092_17969# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X13 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=9.86 ps=87.72 w=1 l=0.4
X14 VOUT VOUT VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X15 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X16 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X17 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X18 VOUT a_6092_17969# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X19 a_6092_17969# VP a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X20 a_6092_17969# VP a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X21 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X22 a_6423_5719# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X23 a_6423_5719# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X24 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X25 a_6105_7756# VN a_6939_14134# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X26 a_6105_7756# VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=1
X27 VOUT VOUT VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X28 VSS a_4943_7756# a_6423_5719# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X29 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X30 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X31 a_6423_5719# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X32 a_6423_5719# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X33 a_6939_14134# VN a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X34 a_6939_14134# VN a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X35 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X36 a_6681_4767# a_7841_7668# VOUT VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X37 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X38 a_6105_7756# VP a_6092_17969# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X39 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X40 VOUT a_6092_17969# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X41 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X42 VOUT EN a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X43 a_6105_7756# VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=1
X44 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X45 VOUT a_6092_17969# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X46 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X47 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X48 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X49 VOUT a_6092_17969# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X50 VDD a_6092_17969# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X51 a_6939_14134# a_6939_14134# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X52 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X53 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X54 VSS a_4943_7756# a_6423_5719# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X55 VDD a_6092_17969# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X56 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X57 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X58 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X59 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X60 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X61 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X62 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X63 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X64 VSS a_4943_7756# a_6423_5719# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X65 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X66 VDD a_6939_14134# a_6092_17969# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X67 a_6423_5719# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X68 VDD a_6939_14134# a_6092_17969# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X69 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X70 a_6939_14134# a_6939_14134# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X71 VOUT a_6092_17969# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X72 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X73 C1 VOUT sky130_fd_pr__cap_mim_m3_1 l=25.5 w=25.5
X74 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X75 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X76 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X77 VSS VSS a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=1
X78 VOUT a_6092_17969# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X79 a_6939_14134# VN a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X80 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X81 IBIAS IBIAS IBIAS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=4.06 ps=29.16 w=7 l=1
X82 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X83 IBIAS EN a_4943_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X84 VOUT a_6092_17969# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X85 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X86 a_6105_7756# VP a_6092_17969# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X87 a_6681_4767# a_6681_4767# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X88 VDD a_6092_17969# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X89 a_4943_7756# a_4943_7756# a_4943_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=4.93 ps=35.74 w=7 l=1
X90 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X91 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X92 VSS VSS a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=1
X93 VDD a_6092_17969# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X94 a_6092_17969# VP a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X95 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X96 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X97 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X98 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X99 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X100 a_6105_7756# VN a_6939_14134# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X101 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X102 VSS a_4943_7756# a_6423_5719# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X103 VSS a_4943_7756# a_6423_5719# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X104 a_6105_7756# VP a_6092_17969# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X105 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X106 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X107 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X108 a_6423_5719# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X109 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X110 VSS a_4943_7756# a_6423_5719# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X111 a_6092_17969# a_6739_12378# a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X112 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X113 VDD a_6092_17969# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X114 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X115 a_6105_7756# VN a_6939_14134# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X116 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X117 VDD a_6092_17969# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X118 a_6105_7756# VN a_6939_14134# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X119 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X120 a_6939_14134# a_6739_14046# a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X121 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X122 VDD a_6092_17969# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X123 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X124 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X125 VOUT VOUT VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X126 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X127 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X128 a_6939_14134# VN a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X129 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X130 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X131 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X132 a_6423_5719# a_6423_5719# a_6423_5719# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=9.28 ps=68.64 w=7 l=1
X133 C1 a_6092_17969# VSS sky130_fd_pr__res_xhigh_po_1p41 l=14
X134 VOUT a_6092_17969# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X135 a_6681_4767# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X136 a_6105_7756# VP a_6092_17969# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X137 VDD a_6939_14134# a_6939_14134# VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X138 a_4943_7756# a_4943_7756# VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X139 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X140 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X141 a_6423_5719# EN a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X142 a_6092_17969# a_6939_14134# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X143 a_6092_17969# a_6939_14134# VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X144 a_6105_7756# a_6105_7756# a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=28.42 ps=204.12 w=7 l=1
X145 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X146 VSS VSS VSS VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X147 a_6105_7756# a_9061_12378# a_6092_17969# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X148 a_6092_17969# VP a_6105_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X149 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X150 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X151 VSS a_4943_7756# a_4943_7756# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X152 VDD a_6092_17969# VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X153 VDD VDD VDD VDD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X154 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X155 VSS a_4943_7756# a_6681_4767# VSS sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
.ends

