* NGSPICE file created from two_stage_op_amp.ext - technology: sky130A

.subckt two_stage_op_amp EN VSS IBIAS VOUT VP VN VDD
X0 a_6681_4767.t26 a_4943_7756.t8 VSS.t122 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X1 VDD.t21 a_6681_14134.t0 a_6681_14134.t1 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X2 VSS.t81 VSS.t80 VSS.t81 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X3 VSS.t79 VSS.t78 VSS.t79 VSS.t68 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X4 VDD.t71 a_6092_17969.t18 VOUT.t28 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X5 VSS.t121 a_4943_7756.t9 a_6681_4767.t25 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 VSS.t77 VSS.t76 VSS.t77 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X7 VSS.t75 VSS.t74 VSS.t75 VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X8 a_6681_4767.t2 a_6681_4767.t0 a_6681_4767.t1 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X9 VOUT.t10 VOUT.t9 VOUT.t10 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X10 a_6681_14134.t8 a_6681_14134.t7 a_6681_14134.t8 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X11 VSS.t73 VSS.t72 VSS.t73 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X12 VOUT.t27 a_6092_17969.t19 VDD.t24 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X13 VDD.t67 VDD.t66 VDD.t67 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X14 VOUT.t8 VOUT.t6 VOUT.t7 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X15 a_6681_4767.t24 a_4943_7756.t10 VSS.t120 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 VSS.t71 VSS.t70 VSS.t71 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X17 VOUT.t26 a_6092_17969.t20 VDD.t76 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X18 a_6092_17969.t16 VP.t0 a_6105_7756.t16 VSS.t68 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X19 a_6092_17969.t10 VP.t1 a_6105_7756.t15 VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X20 a_6681_4767.t23 a_4943_7756.t11 VSS.t119 VSS.t106 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X21 a_6423_5719.t13 a_4943_7756.t12 VSS.t118 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X22 a_6423_5719.t12 a_4943_7756.t13 VSS.t117 VSS.t68 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X23 VSS.t116 a_4943_7756.t14 a_6681_4767.t22 VSS.t103 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X24 a_6105_7756.t3 VN.t0 a_6681_14134.t13 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X25 VOUT.t5 VOUT.t4 VOUT.t5 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X26 VSS.t115 a_4943_7756.t15 a_6423_5719.t11 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X27 VDD.t65 VDD.t63 VDD.t64 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X28 a_6681_4767.t21 a_4943_7756.t16 VSS.t114 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X29 a_6423_5719.t10 a_4943_7756.t17 VSS.t113 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X30 a_6423_5719.t9 a_4943_7756.t18 VSS.t112 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X31 a_6681_14134.t20 VN.t1 a_6105_7756.t19 VSS.t68 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X32 a_6681_14134.t14 VN.t2 a_6105_7756.t4 VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X33 VOUT.t3 VOUT.t2 VOUT.t3 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X34 VSS.t69 VSS.t67 VSS.t69 VSS.t68 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X35 a_6681_4767.t20 a_4943_7756.t19 VSS.t111 VSS.t106 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X36 a_6105_7756.t14 VP.t2 a_6092_17969.t12 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X37 VSS.t66 VSS.t64 VSS.t66 VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X38 VOUT.t25 a_6092_17969.t21 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X39 VSS.t110 a_4943_7756.t20 a_6681_4767.t19 VSS.t103 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X40 VOUT.t30 EN.t0 a_6681_4767.t27 VSS.t127 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X41 VDD.t62 VDD.t60 VDD.t61 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X42 VOUT.t24 a_6092_17969.t22 VDD.t73 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X43 VSS.t63 VSS.t61 VSS.t63 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X44 VDD.t59 VDD.t58 VDD.t59 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X45 VOUT.t23 a_6092_17969.t23 VDD.t74 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X46 VDD.t75 a_6092_17969.t24 VOUT.t22 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X47 a_6681_14134.t10 a_6681_14134.t9 VDD.t20 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X48 VSS.t60 VSS.t59 VSS.t60 VSS.t35 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X49 VDD.t57 VDD.t56 VDD.t57 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X50 VSS.t109 a_4943_7756.t21 a_6423_5719.t8 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X51 VDD.t8 a_6092_17969.t25 VOUT.t21 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X52 VSS.t58 VSS.t57 VSS.t58 VSS.t49 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X53 a_6681_4767.t18 a_4943_7756.t22 VSS.t108 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X54 VDD.t55 VDD.t54 VDD.t55 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X55 VDD.t53 VDD.t52 VDD.t53 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X56 VSS.t102 a_4943_7756.t23 a_6681_4767.t17 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X57 VSS.t56 VSS.t55 VSS.t56 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X58 VDD.t51 VDD.t50 VDD.t51 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X59 VSS.t107 a_4943_7756.t24 a_6423_5719.t7 VSS.t106 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X60 a_6681_4767.t16 a_4943_7756.t25 VSS.t105 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X61 VDD.t19 a_6681_14134.t21 a_6092_17969.t3 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X62 a_6423_5719.t6 a_4943_7756.t26 VSS.t104 VSS.t103 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X63 VDD.t18 a_6681_14134.t22 a_6092_17969.t2 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X64 VSS.t54 VSS.t53 VSS.t54 VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X65 a_6681_14134.t3 a_6681_14134.t2 VDD.t16 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X66 VOUT.t20 a_6092_17969.t26 VDD.t9 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X67 VSS.t52 VSS.t51 VSS.t52 VSS.t35 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X68 C1.t1 VOUT.t29 sky130_fd_pr__cap_mim_m3_1 l=25.5 w=25.5
X69 VSS.t50 VSS.t48 VSS.t50 VSS.t49 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X70 VDD.t49 VDD.t48 VDD.t49 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X71 a_6681_4767.t15 a_4943_7756.t27 VSS.t101 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X72 VOUT.t19 a_6092_17969.t27 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X73 a_6681_14134.t16 VN.t3 a_6105_7756.t6 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X74 VSS.t100 a_4943_7756.t28 a_6681_4767.t14 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X75 IBIAS.t2 IBIAS.t1 IBIAS.t2 VSS.t128 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X76 VDD.t47 VDD.t46 VDD.t47 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X77 IBIAS.t0 EN.t1 a_4943_7756.t7 VSS.t125 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X78 VOUT.t18 a_6092_17969.t28 VDD.t72 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X79 a_6681_4767.t13 a_4943_7756.t29 VSS.t99 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X80 a_6105_7756.t13 VP.t3 a_6092_17969.t13 VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X81 VDD.t1 a_6092_17969.t29 VOUT.t17 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X82 a_4943_7756.t2 a_4943_7756.t0 a_4943_7756.t1 VSS.t98 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X83 VSS.t47 VSS.t46 VSS.t47 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X84 VSS.t45 VSS.t43 VSS.t44 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X85 VDD.t10 a_6092_17969.t30 VOUT.t16 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X86 a_6092_17969.t14 VP.t4 a_6105_7756.t12 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X87 VSS.t97 a_4943_7756.t30 a_6681_4767.t12 VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X88 VSS.t42 VSS.t40 VSS.t41 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X89 VDD.t45 VDD.t42 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X90 a_6105_7756.t7 VN.t4 a_6681_14134.t17 VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X91 VSS.t39 VSS.t37 VSS.t39 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X92 VSS.t36 VSS.t34 VSS.t36 VSS.t35 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X93 VSS.t94 a_4943_7756.t31 a_6423_5719.t5 VSS.t49 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X94 VSS.t96 a_4943_7756.t32 a_6423_5719.t4 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X95 a_6105_7756.t11 VP.t5 a_6092_17969.t15 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X96 a_6681_4767.t11 a_4943_7756.t33 VSS.t95 VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X97 VSS.t33 VSS.t31 VSS.t32 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X98 a_6423_5719.t3 a_4943_7756.t34 VSS.t93 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X99 VSS.t30 VSS.t28 VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X100 VSS.t27 VSS.t26 VSS.t27 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X101 VSS.t92 a_4943_7756.t35 a_6423_5719.t2 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X102 a_6092_17969.t9 a_6092_17969.t7 a_6092_17969.t8 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X103 VSS.t91 a_4943_7756.t36 a_6681_4767.t10 VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X104 VDD.t68 a_6092_17969.t31 VOUT.t15 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X105 VSS.t25 VSS.t24 VSS.t25 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X106 a_6105_7756.t18 VN.t5 a_6681_14134.t19 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X107 a_6681_4767.t9 a_4943_7756.t37 VSS.t90 VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X108 VDD.t25 a_6092_17969.t32 VOUT.t14 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X109 a_6105_7756.t17 VN.t6 a_6681_14134.t18 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X110 VSS.t23 VSS.t21 VSS.t23 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X111 a_6681_14134.t6 a_6681_14134.t4 a_6681_14134.t5 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X112 VDD.t41 VDD.t40 VDD.t41 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X113 VDD.t69 a_6092_17969.t33 VOUT.t13 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X114 VSS.t20 VSS.t18 VSS.t20 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X115 VDD.t39 VDD.t38 VDD.t39 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X116 VOUT.t1 VOUT.t0 VOUT.t1 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X117 VSS.t17 VSS.t15 VSS.t16 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X118 VSS.t89 a_4943_7756.t38 a_6681_4767.t8 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X119 a_6681_14134.t15 VN.t7 a_6105_7756.t5 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X120 VDD.t37 VDD.t36 VDD.t37 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X121 VSS.t88 a_4943_7756.t39 a_6681_4767.t7 VSS.t68 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X122 VSS.t14 VSS.t11 VSS.t13 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X123 a_6423_5719.t1 a_6423_5719.t0 a_6423_5719.t1 VSS.t124 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X124 C1.t0 a_6092_17969.t11 VSS.t123 sky130_fd_pr__res_xhigh_po_1p41 l=14
X125 VOUT.t12 a_6092_17969.t34 VDD.t70 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X126 a_6681_4767.t6 a_4943_7756.t40 VSS.t86 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X127 a_6105_7756.t10 VP.t6 a_6092_17969.t17 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X128 VDD.t15 a_6681_14134.t11 a_6681_14134.t12 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X129 a_4943_7756.t6 a_4943_7756.t5 VSS.t87 VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X130 VSS.t85 a_4943_7756.t41 a_6681_4767.t5 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X131 VSS.t10 VSS.t8 VSS.t10 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X132 a_6423_5719.t14 EN.t2 a_6105_7756.t8 VSS.t126 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X133 a_6092_17969.t1 a_6681_14134.t23 VDD.t13 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X134 a_6092_17969.t0 a_6681_14134.t24 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X135 a_6105_7756.t2 a_6105_7756.t0 a_6105_7756.t1 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X136 VDD.t35 VDD.t33 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X137 VSS.t7 VSS.t5 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X138 a_6092_17969.t6 a_6092_17969.t5 a_6092_17969.t6 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X139 a_6092_17969.t4 VP.t7 a_6105_7756.t9 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X140 VDD.t32 VDD.t31 VDD.t32 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X141 VDD.t30 VDD.t28 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X142 VSS.t83 a_4943_7756.t3 a_4943_7756.t4 VSS.t29 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X143 VDD.t23 a_6092_17969.t35 VOUT.t11 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X144 VDD.t27 VDD.t26 VDD.t27 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X145 VSS.t84 a_4943_7756.t42 a_6681_4767.t4 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X146 VSS.t82 a_4943_7756.t43 a_6681_4767.t3 VSS.t68 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
C0 EN IBIAS 0.80215f
C1 C1 VOUT 57.5804f
C2 VP VOUT 0.11738f
C3 EN VOUT 0.50424f
C4 VP VN 5.95617f
C5 VDD VOUT 9.39455f
R0 a_4943_7756.n87 a_4943_7756.n86 185
R1 a_4943_7756.n86 a_4943_7756.n85 185
R2 a_4943_7756.n86 a_4943_7756.n8 185
R3 a_4943_7756.n86 a_4943_7756.n7 185
R4 a_4943_7756.n86 a_4943_7756.n6 185
R5 a_4943_7756.n86 a_4943_7756.n5 185
R6 a_4943_7756.n86 a_4943_7756.n4 185
R7 a_4943_7756.n42 a_4943_7756.n41 185
R8 a_4943_7756.n42 a_4943_7756.n29 185
R9 a_4943_7756.n42 a_4943_7756.n28 185
R10 a_4943_7756.n42 a_4943_7756.n26 185
R11 a_4943_7756.n42 a_4943_7756.n25 185
R12 a_4943_7756.n43 a_4943_7756.n42 185
R13 a_4943_7756.t2 a_4943_7756.n92 180.167
R14 a_4943_7756.t2 a_4943_7756.n92 180.167
R15 a_4943_7756.n60 a_4943_7756.t20 165.607
R16 a_4943_7756.n10 a_4943_7756.t31 165.607
R17 a_4943_7756.n70 a_4943_7756.t19 165.032
R18 a_4943_7756.n69 a_4943_7756.t42 165.032
R19 a_4943_7756.n68 a_4943_7756.t16 165.032
R20 a_4943_7756.n67 a_4943_7756.t28 165.032
R21 a_4943_7756.n66 a_4943_7756.t27 165.032
R22 a_4943_7756.n65 a_4943_7756.t36 165.032
R23 a_4943_7756.n64 a_4943_7756.t37 165.032
R24 a_4943_7756.n63 a_4943_7756.t9 165.032
R25 a_4943_7756.n62 a_4943_7756.t8 165.032
R26 a_4943_7756.n61 a_4943_7756.t43 165.032
R27 a_4943_7756.n60 a_4943_7756.t29 165.032
R28 a_4943_7756.n59 a_4943_7756.t18 165.032
R29 a_4943_7756.n57 a_4943_7756.t11 163.058
R30 a_4943_7756.n55 a_4943_7756.t38 163.058
R31 a_4943_7756.n53 a_4943_7756.t10 163.058
R32 a_4943_7756.n51 a_4943_7756.t23 163.058
R33 a_4943_7756.n49 a_4943_7756.t22 163.058
R34 a_4943_7756.n21 a_4943_7756.t33 163.058
R35 a_4943_7756.n47 a_4943_7756.t30 163.058
R36 a_4943_7756.n17 a_4943_7756.t41 163.058
R37 a_4943_7756.n15 a_4943_7756.t40 163.058
R38 a_4943_7756.n13 a_4943_7756.t39 163.058
R39 a_4943_7756.n11 a_4943_7756.t25 163.058
R40 a_4943_7756.n9 a_4943_7756.t14 163.058
R41 a_4943_7756.t5 a_4943_7756.n45 162.941
R42 a_4943_7756.n45 a_4943_7756.t3 162.941
R43 a_4943_7756.n57 a_4943_7756.t24 162.781
R44 a_4943_7756.n55 a_4943_7756.t12 162.781
R45 a_4943_7756.n53 a_4943_7756.t21 162.781
R46 a_4943_7756.n51 a_4943_7756.t34 162.781
R47 a_4943_7756.n49 a_4943_7756.t32 162.781
R48 a_4943_7756.n17 a_4943_7756.t17 162.781
R49 a_4943_7756.n15 a_4943_7756.t15 162.781
R50 a_4943_7756.n13 a_4943_7756.t13 162.781
R51 a_4943_7756.n11 a_4943_7756.t35 162.781
R52 a_4943_7756.n9 a_4943_7756.t26 162.781
R53 a_4943_7756.n46 a_4943_7756.t5 162.639
R54 a_4943_7756.t3 a_4943_7756.n22 162.639
R55 a_4943_7756.n91 a_4943_7756.t0 130.75
R56 a_4943_7756.n86 a_4943_7756.n3 86.5152
R57 a_4943_7756.n42 a_4943_7756.n27 86.5152
R58 a_4943_7756.n88 a_4943_7756.n0 30.3012
R59 a_4943_7756.n73 a_4943_7756.n4 24.8476
R60 a_4943_7756.n35 a_4943_7756.n28 24.8476
R61 a_4943_7756.n33 a_4943_7756.n26 24.8476
R62 a_4943_7756.n75 a_4943_7756.n5 23.3417
R63 a_4943_7756.n37 a_4943_7756.n29 23.3417
R64 a_4943_7756.n31 a_4943_7756.n25 23.3417
R65 a_4943_7756.n72 a_4943_7756.n3 22.0256
R66 a_4943_7756.n77 a_4943_7756.n6 21.8358
R67 a_4943_7756.n41 a_4943_7756.n40 21.8358
R68 a_4943_7756.n43 a_4943_7756.n24 21.8358
R69 a_4943_7756.n79 a_4943_7756.n7 20.3299
R70 a_4943_7756.n81 a_4943_7756.n8 18.824
R71 a_4943_7756.n85 a_4943_7756.n84 17.3181
R72 a_4943_7756.n86 a_4943_7756.n0 16.3559
R73 a_4943_7756.n87 a_4943_7756.n2 15.8123
R74 a_4943_7756.n41 a_4943_7756.n30 14.5711
R75 a_4943_7756.n44 a_4943_7756.n43 14.5711
R76 a_4943_7756.n73 a_4943_7756.n3 12.7256
R77 a_4943_7756.n35 a_4943_7756.n27 12.7256
R78 a_4943_7756.n33 a_4943_7756.n27 12.7256
R79 a_4943_7756.n88 a_4943_7756.n87 11.2946
R80 a_4943_7756.n85 a_4943_7756.n2 9.78874
R81 a_4943_7756.n36 a_4943_7756.n35 9.3005
R82 a_4943_7756.n38 a_4943_7756.n37 9.3005
R83 a_4943_7756.n40 a_4943_7756.n39 9.3005
R84 a_4943_7756.n34 a_4943_7756.n33 9.3005
R85 a_4943_7756.n32 a_4943_7756.n31 9.3005
R86 a_4943_7756.n24 a_4943_7756.n23 9.3005
R87 a_4943_7756.n74 a_4943_7756.n73 9.3005
R88 a_4943_7756.n76 a_4943_7756.n75 9.3005
R89 a_4943_7756.n78 a_4943_7756.n77 9.3005
R90 a_4943_7756.n80 a_4943_7756.n79 9.3005
R91 a_4943_7756.n82 a_4943_7756.n81 9.3005
R92 a_4943_7756.n84 a_4943_7756.n83 9.3005
R93 a_4943_7756.n2 a_4943_7756.n1 9.3005
R94 a_4943_7756.n89 a_4943_7756.n88 9.3005
R95 a_4943_7756.n84 a_4943_7756.n8 8.28285
R96 a_4943_7756.n81 a_4943_7756.n7 6.77697
R97 a_4943_7756.n42 a_4943_7756.t4 5.8005
R98 a_4943_7756.n42 a_4943_7756.t6 5.8005
R99 a_4943_7756.n71 a_4943_7756.n70 5.72243
R100 a_4943_7756.n79 a_4943_7756.n6 5.27109
R101 a_4943_7756.n72 a_4943_7756.n71 4.70369
R102 a_4943_7756.n71 a_4943_7756.n59 4.58132
R103 a_4943_7756.n77 a_4943_7756.n5 3.76521
R104 a_4943_7756.n40 a_4943_7756.n29 3.76521
R105 a_4943_7756.n25 a_4943_7756.n24 3.76521
R106 a_4943_7756.n86 a_4943_7756.t7 2.48621
R107 a_4943_7756.n86 a_4943_7756.t1 2.48621
R108 a_4943_7756.n90 a_4943_7756.n0 2.36936
R109 a_4943_7756.n75 a_4943_7756.n4 2.25932
R110 a_4943_7756.n37 a_4943_7756.n28 2.25932
R111 a_4943_7756.n31 a_4943_7756.n26 2.25932
R112 a_4943_7756.n58 a_4943_7756.n57 2.25162
R113 a_4943_7756.n56 a_4943_7756.n55 2.25162
R114 a_4943_7756.n54 a_4943_7756.n53 2.25162
R115 a_4943_7756.n52 a_4943_7756.n51 2.25162
R116 a_4943_7756.n50 a_4943_7756.n49 2.25162
R117 a_4943_7756.n21 a_4943_7756.n19 2.25162
R118 a_4943_7756.n48 a_4943_7756.n47 2.25162
R119 a_4943_7756.n18 a_4943_7756.n17 2.25162
R120 a_4943_7756.n16 a_4943_7756.n15 2.25162
R121 a_4943_7756.n14 a_4943_7756.n13 2.25162
R122 a_4943_7756.n12 a_4943_7756.n11 2.25162
R123 a_4943_7756.n10 a_4943_7756.n9 2.25162
R124 a_4943_7756.n92 a_4943_7756.n91 1.27148
R125 a_4943_7756.n61 a_4943_7756.n60 0.574917
R126 a_4943_7756.n62 a_4943_7756.n61 0.574917
R127 a_4943_7756.n63 a_4943_7756.n62 0.574917
R128 a_4943_7756.n64 a_4943_7756.n63 0.574917
R129 a_4943_7756.n65 a_4943_7756.n64 0.574917
R130 a_4943_7756.n66 a_4943_7756.n65 0.574917
R131 a_4943_7756.n67 a_4943_7756.n66 0.574917
R132 a_4943_7756.n68 a_4943_7756.n67 0.574917
R133 a_4943_7756.n69 a_4943_7756.n68 0.574917
R134 a_4943_7756.n70 a_4943_7756.n69 0.574917
R135 a_4943_7756.n12 a_4943_7756.n10 0.574917
R136 a_4943_7756.n14 a_4943_7756.n12 0.574917
R137 a_4943_7756.n16 a_4943_7756.n14 0.574917
R138 a_4943_7756.n18 a_4943_7756.n16 0.574917
R139 a_4943_7756.n19 a_4943_7756.n18 0.574917
R140 a_4943_7756.n48 a_4943_7756.n19 0.574917
R141 a_4943_7756.n50 a_4943_7756.n48 0.574917
R142 a_4943_7756.n52 a_4943_7756.n50 0.574917
R143 a_4943_7756.n54 a_4943_7756.n52 0.574917
R144 a_4943_7756.n56 a_4943_7756.n54 0.574917
R145 a_4943_7756.n58 a_4943_7756.n56 0.574917
R146 a_4943_7756.n59 a_4943_7756.n58 0.574917
R147 a_4943_7756.n91 a_4943_7756.n90 0.320353
R148 a_4943_7756.n22 a_4943_7756.n20 0.302413
R149 a_4943_7756.n46 a_4943_7756.n20 0.302413
R150 a_4943_7756.n30 a_4943_7756.n20 0.217891
R151 a_4943_7756.n45 a_4943_7756.n44 0.217891
R152 a_4943_7756.n39 a_4943_7756.n30 0.196152
R153 a_4943_7756.n39 a_4943_7756.n38 0.196152
R154 a_4943_7756.n38 a_4943_7756.n36 0.196152
R155 a_4943_7756.n36 a_4943_7756.n34 0.196152
R156 a_4943_7756.n34 a_4943_7756.n32 0.196152
R157 a_4943_7756.n32 a_4943_7756.n23 0.196152
R158 a_4943_7756.n44 a_4943_7756.n23 0.196152
R159 a_4943_7756.n90 a_4943_7756.n89 0.196152
R160 a_4943_7756.n89 a_4943_7756.n1 0.196152
R161 a_4943_7756.n83 a_4943_7756.n1 0.196152
R162 a_4943_7756.n83 a_4943_7756.n82 0.196152
R163 a_4943_7756.n82 a_4943_7756.n80 0.196152
R164 a_4943_7756.n80 a_4943_7756.n78 0.196152
R165 a_4943_7756.n78 a_4943_7756.n76 0.196152
R166 a_4943_7756.n76 a_4943_7756.n74 0.196152
R167 a_4943_7756.n74 a_4943_7756.n72 0.196152
R168 a_4943_7756.n22 a_4943_7756.n21 0.142018
R169 a_4943_7756.n47 a_4943_7756.n46 0.142018
R170 VSS.n1049 VSS.n305 4887.33
R171 VSS.n248 VSS.n236 1321.06
R172 VSS.n2248 VSS.n2159 1321.06
R173 VSS.n2315 VSS.n2314 1321.06
R174 VSS.n245 VSS.n234 1321.06
R175 VSS.n2142 VSS.n564 1268.91
R176 VSS.n2117 VSS.n582 1268.91
R177 VSS.n652 VSS.n562 1268.91
R178 VSS.n2074 VSS.n584 1268.91
R179 VSS.n1726 VSS.n810 1268.91
R180 VSS.n2296 VSS.n339 1268.91
R181 VSS.n1779 VSS.n1714 1268.91
R182 VSS.n2253 VSS.n2252 1268.91
R183 VSS.n1635 VSS.n957 1268.91
R184 VSS.n2052 VSS.n737 1268.91
R185 VSS.n1592 VSS.n1591 1268.91
R186 VSS.n2054 VSS.n733 1268.91
R187 VSS.n1148 VSS.n1051 1182
R188 VSS.n2150 VSS.n368 1182
R189 VSS.n1073 VSS.n1047 1182
R190 VSS.n2152 VSS.n366 1182
R191 VSS.n1232 VSS.n1018 1182
R192 VSS.n1989 VSS.n889 1182
R193 VSS.n1803 VSS.n886 1182
R194 VSS.n1429 VSS.n1028 1182
R195 VSS.n1946 VSS.n1945 996.588
R196 VSS.n1898 VSS.n1897 602.588
R197 VSS.n1850 VSS.n1849 602.588
R198 VSS.n245 VSS.n244 585
R199 VSS.n246 VSS.n245 585
R200 VSS.n243 VSS.n240 585
R201 VSS.n242 VSS.n241 585
R202 VSS.n238 VSS.n237 585
R203 VSS.n249 VSS.n248 585
R204 VSS.n2368 VSS.n2367 585
R205 VSS.n2369 VSS.n2368 585
R206 VSS.n301 VSS.n300 585
R207 VSS.n2370 VSS.n301 585
R208 VSS.n2373 VSS.n2372 585
R209 VSS.n2372 VSS.n2371 585
R210 VSS.n2374 VSS.n299 585
R211 VSS.n299 VSS.n298 585
R212 VSS.n2376 VSS.n2375 585
R213 VSS.n2377 VSS.n2376 585
R214 VSS.n294 VSS.n293 585
R215 VSS.n2378 VSS.n294 585
R216 VSS.n2381 VSS.n2380 585
R217 VSS.n2380 VSS.n2379 585
R218 VSS.n2382 VSS.n208 585
R219 VSS.n208 VSS.n206 585
R220 VSS.n2384 VSS.n2383 585
R221 VSS.n2385 VSS.n2384 585
R222 VSS.n292 VSS.n207 585
R223 VSS.n207 VSS.n205 585
R224 VSS.n291 VSS.n290 585
R225 VSS.n290 VSS.n289 585
R226 VSS.n210 VSS.n209 585
R227 VSS.n211 VSS.n210 585
R228 VSS.n282 VSS.n281 585
R229 VSS.n283 VSS.n282 585
R230 VSS.n280 VSS.n216 585
R231 VSS.n216 VSS.n215 585
R232 VSS.n279 VSS.n278 585
R233 VSS.n278 VSS.n277 585
R234 VSS.n218 VSS.n217 585
R235 VSS.n219 VSS.n218 585
R236 VSS.n270 VSS.n269 585
R237 VSS.n271 VSS.n270 585
R238 VSS.n268 VSS.n224 585
R239 VSS.n224 VSS.n223 585
R240 VSS.n267 VSS.n266 585
R241 VSS.n266 VSS.n265 585
R242 VSS.n226 VSS.n225 585
R243 VSS.n227 VSS.n226 585
R244 VSS.n258 VSS.n257 585
R245 VSS.n259 VSS.n258 585
R246 VSS.n256 VSS.n232 585
R247 VSS.n232 VSS.n231 585
R248 VSS.n255 VSS.n254 585
R249 VSS.n254 VSS.n253 585
R250 VSS.n234 VSS.n233 585
R251 VSS.n235 VSS.n234 585
R252 VSS.n250 VSS.n236 585
R253 VSS.n236 VSS.n235 585
R254 VSS.n252 VSS.n251 585
R255 VSS.n253 VSS.n252 585
R256 VSS.n230 VSS.n229 585
R257 VSS.n231 VSS.n230 585
R258 VSS.n261 VSS.n260 585
R259 VSS.n260 VSS.n259 585
R260 VSS.n262 VSS.n228 585
R261 VSS.n228 VSS.n227 585
R262 VSS.n264 VSS.n263 585
R263 VSS.n265 VSS.n264 585
R264 VSS.n222 VSS.n221 585
R265 VSS.n223 VSS.n222 585
R266 VSS.n273 VSS.n272 585
R267 VSS.n272 VSS.n271 585
R268 VSS.n274 VSS.n220 585
R269 VSS.n220 VSS.n219 585
R270 VSS.n276 VSS.n275 585
R271 VSS.n277 VSS.n276 585
R272 VSS.n214 VSS.n213 585
R273 VSS.n215 VSS.n214 585
R274 VSS.n285 VSS.n284 585
R275 VSS.n284 VSS.n283 585
R276 VSS.n286 VSS.n212 585
R277 VSS.n212 VSS.n211 585
R278 VSS.n288 VSS.n287 585
R279 VSS.n289 VSS.n288 585
R280 VSS.n203 VSS.n201 585
R281 VSS.n205 VSS.n203 585
R282 VSS.n2387 VSS.n2386 585
R283 VSS.n2386 VSS.n2385 585
R284 VSS.n204 VSS.n202 585
R285 VSS.n206 VSS.n204 585
R286 VSS.n2181 VSS.n295 585
R287 VSS.n2379 VSS.n295 585
R288 VSS.n2182 VSS.n296 585
R289 VSS.n2378 VSS.n296 585
R290 VSS.n2183 VSS.n297 585
R291 VSS.n2377 VSS.n297 585
R292 VSS.n2185 VSS.n2184 585
R293 VSS.n2184 VSS.n298 585
R294 VSS.n2186 VSS.n302 585
R295 VSS.n2371 VSS.n302 585
R296 VSS.n2187 VSS.n303 585
R297 VSS.n2370 VSS.n303 585
R298 VSS.n2188 VSS.n304 585
R299 VSS.n2369 VSS.n304 585
R300 VSS.n2240 VSS.n2239 585
R301 VSS.n2238 VSS.n2180 585
R302 VSS.n2237 VSS.n2179 585
R303 VSS.n2242 VSS.n2179 585
R304 VSS.n2236 VSS.n2235 585
R305 VSS.n2234 VSS.n2233 585
R306 VSS.n2232 VSS.n2231 585
R307 VSS.n2230 VSS.n2229 585
R308 VSS.n2228 VSS.n2227 585
R309 VSS.n2226 VSS.n2225 585
R310 VSS.n2224 VSS.n2223 585
R311 VSS.n2222 VSS.n2221 585
R312 VSS.n2220 VSS.n2219 585
R313 VSS.n2218 VSS.n2217 585
R314 VSS.n2216 VSS.n2215 585
R315 VSS.n2214 VSS.n2213 585
R316 VSS.n2212 VSS.n2211 585
R317 VSS.n2210 VSS.n2209 585
R318 VSS.n2208 VSS.n2207 585
R319 VSS.n2206 VSS.n2205 585
R320 VSS.n2204 VSS.n2203 585
R321 VSS.n2202 VSS.n2201 585
R322 VSS.n2200 VSS.n2199 585
R323 VSS.n2198 VSS.n2197 585
R324 VSS.n2196 VSS.n2195 585
R325 VSS.n2194 VSS.n2193 585
R326 VSS.n2192 VSS.n2191 585
R327 VSS.n2190 VSS.n2189 585
R328 VSS.n2165 VSS.n2164 585
R329 VSS.n2245 VSS.n2244 585
R330 VSS.n2246 VSS.n2159 585
R331 VSS.n2242 VSS.n2159 585
R332 VSS.n2316 VSS.n2315 585
R333 VSS.n2317 VSS.n328 585
R334 VSS.n2319 VSS.n2318 585
R335 VSS.n2321 VSS.n326 585
R336 VSS.n2323 VSS.n2322 585
R337 VSS.n2324 VSS.n325 585
R338 VSS.n2326 VSS.n2325 585
R339 VSS.n2328 VSS.n323 585
R340 VSS.n2330 VSS.n2329 585
R341 VSS.n2331 VSS.n322 585
R342 VSS.n2333 VSS.n2332 585
R343 VSS.n2335 VSS.n320 585
R344 VSS.n2337 VSS.n2336 585
R345 VSS.n2338 VSS.n319 585
R346 VSS.n2340 VSS.n2339 585
R347 VSS.n2342 VSS.n317 585
R348 VSS.n2344 VSS.n2343 585
R349 VSS.n2345 VSS.n316 585
R350 VSS.n2347 VSS.n2346 585
R351 VSS.n2349 VSS.n314 585
R352 VSS.n2351 VSS.n2350 585
R353 VSS.n2352 VSS.n313 585
R354 VSS.n2354 VSS.n2353 585
R355 VSS.n2356 VSS.n311 585
R356 VSS.n2358 VSS.n2357 585
R357 VSS.n2359 VSS.n310 585
R358 VSS.n2361 VSS.n2360 585
R359 VSS.n2363 VSS.n307 585
R360 VSS.n2365 VSS.n2364 585
R361 VSS.n2366 VSS.n306 585
R362 VSS.n2148 VSS.n368 585
R363 VSS.n2147 VSS.n2146 585
R364 VSS.n370 VSS.n369 585
R365 VSS.n2144 VSS.n370 585
R366 VSS.n391 VSS.n390 585
R367 VSS.n393 VSS.n392 585
R368 VSS.n395 VSS.n394 585
R369 VSS.n397 VSS.n396 585
R370 VSS.n399 VSS.n398 585
R371 VSS.n401 VSS.n400 585
R372 VSS.n403 VSS.n402 585
R373 VSS.n405 VSS.n404 585
R374 VSS.n407 VSS.n406 585
R375 VSS.n409 VSS.n408 585
R376 VSS.n411 VSS.n410 585
R377 VSS.n413 VSS.n412 585
R378 VSS.n415 VSS.n414 585
R379 VSS.n417 VSS.n416 585
R380 VSS.n419 VSS.n418 585
R381 VSS.n421 VSS.n420 585
R382 VSS.n423 VSS.n422 585
R383 VSS.n425 VSS.n424 585
R384 VSS.n427 VSS.n426 585
R385 VSS.n430 VSS.n429 585
R386 VSS.n428 VSS.n389 585
R387 VSS.n534 VSS.n533 585
R388 VSS.n536 VSS.n535 585
R389 VSS.n538 VSS.n537 585
R390 VSS.n540 VSS.n539 585
R391 VSS.n542 VSS.n541 585
R392 VSS.n544 VSS.n543 585
R393 VSS.n546 VSS.n545 585
R394 VSS.n548 VSS.n547 585
R395 VSS.n550 VSS.n549 585
R396 VSS.n552 VSS.n551 585
R397 VSS.n554 VSS.n553 585
R398 VSS.n556 VSS.n555 585
R399 VSS.n557 VSS.n388 585
R400 VSS.n560 VSS.n559 585
R401 VSS.n558 VSS.n366 585
R402 VSS.n2152 VSS.n365 585
R403 VSS.n2152 VSS.n2151 585
R404 VSS.n2154 VSS.n2153 585
R405 VSS.n2153 VSS.n360 585
R406 VSS.n2155 VSS.n349 585
R407 VSS.n2299 VSS.n349 585
R408 VSS.n2157 VSS.n2156 585
R409 VSS.n2250 VSS.n2157 585
R410 VSS.n364 VSS.n342 585
R411 VSS.n2305 VSS.n342 585
R412 VSS.n2001 VSS.n2000 585
R413 VSS.n2002 VSS.n2001 585
R414 VSS.n1999 VSS.n839 585
R415 VSS.n839 VSS.n334 585
R416 VSS.n1998 VSS.n1997 585
R417 VSS.n1997 VSS.n332 585
R418 VSS.n1996 VSS.n835 585
R419 VSS.n2012 VSS.n835 585
R420 VSS.n1995 VSS.n833 585
R421 VSS.n2018 VSS.n833 585
R422 VSS.n1994 VSS.n1993 585
R423 VSS.n1993 VSS.n1992 585
R424 VSS.n840 VSS.n817 585
R425 VSS.n2024 VSS.n817 585
R426 VSS.n1798 VSS.n1797 585
R427 VSS.n1799 VSS.n1798 585
R428 VSS.n1796 VSS.n893 585
R429 VSS.n893 VSS.n809 585
R430 VSS.n1795 VSS.n1794 585
R431 VSS.n1794 VSS.n806 585
R432 VSS.n1793 VSS.n1792 585
R433 VSS.n1793 VSS.n800 585
R434 VSS.n1791 VSS.n798 585
R435 VSS.n2039 VSS.n798 585
R436 VSS.n1790 VSS.n1789 585
R437 VSS.n1789 VSS.n1788 585
R438 VSS.n894 VSS.n790 585
R439 VSS.n2045 VSS.n790 585
R440 VSS.n1452 VSS.n1451 585
R441 VSS.n1452 VSS.n898 585
R442 VSS.n1454 VSS.n1453 585
R443 VSS.n1453 VSS.n735 585
R444 VSS.n1455 VSS.n905 585
R445 VSS.n1697 VSS.n905 585
R446 VSS.n1457 VSS.n1456 585
R447 VSS.n1456 VSS.n903 585
R448 VSS.n1458 VSS.n911 585
R449 VSS.n1690 VSS.n911 585
R450 VSS.n1459 VSS.n920 585
R451 VSS.n1681 VSS.n920 585
R452 VSS.n1460 VSS.n927 585
R453 VSS.n1672 VSS.n927 585
R454 VSS.n1462 VSS.n1461 585
R455 VSS.n1461 VSS.n935 585
R456 VSS.n1463 VSS.n932 585
R457 VSS.n1666 VSS.n932 585
R458 VSS.n1464 VSS.n941 585
R459 VSS.n1657 VSS.n941 585
R460 VSS.n1465 VSS.n948 585
R461 VSS.n1648 VSS.n948 585
R462 VSS.n1467 VSS.n1466 585
R463 VSS.n1466 VSS.n956 585
R464 VSS.n1468 VSS.n953 585
R465 VSS.n1642 VSS.n953 585
R466 VSS.n1470 VSS.n1469 585
R467 VSS.n1469 VSS.n974 585
R468 VSS.n1471 VSS.n961 585
R469 VSS.n1568 VSS.n961 585
R470 VSS.n1473 VSS.n1472 585
R471 VSS.n1472 VSS.n969 585
R472 VSS.n1474 VSS.n967 585
R473 VSS.n1562 VSS.n967 585
R474 VSS.n1477 VSS.n1475 585
R475 VSS.n1477 VSS.n1476 585
R476 VSS.n1479 VSS.n1478 585
R477 VSS.n1478 VSS.n978 585
R478 VSS.n1480 VSS.n984 585
R479 VSS.n1524 VSS.n984 585
R480 VSS.n1482 VSS.n1481 585
R481 VSS.n1481 VSS.n982 585
R482 VSS.n1483 VSS.n991 585
R483 VSS.n1517 VSS.n991 585
R484 VSS.n1485 VSS.n1484 585
R485 VSS.n1485 VSS.n996 585
R486 VSS.n1487 VSS.n1486 585
R487 VSS.n1486 VSS.n995 585
R488 VSS.n1488 VSS.n1002 585
R489 VSS.n1500 VSS.n1002 585
R490 VSS.n1490 VSS.n1489 585
R491 VSS.n1491 VSS.n1490 585
R492 VSS.n1450 VSS.n1009 585
R493 VSS.n1493 VSS.n1009 585
R494 VSS.n1449 VSS.n1448 585
R495 VSS.n1448 VSS.n1447 585
R496 VSS.n1012 VSS.n1011 585
R497 VSS.n1013 VSS.n1012 585
R498 VSS.n1169 VSS.n1021 585
R499 VSS.n1438 VSS.n1021 585
R500 VSS.n1171 VSS.n1170 585
R501 VSS.n1170 VSS.n1019 585
R502 VSS.n1172 VSS.n1027 585
R503 VSS.n1431 VSS.n1027 585
R504 VSS.n1174 VSS.n1173 585
R505 VSS.n1173 VSS.n1026 585
R506 VSS.n1175 VSS.n1032 585
R507 VSS.n1185 VSS.n1032 585
R508 VSS.n1176 VSS.n1038 585
R509 VSS.n1038 VSS.n1031 585
R510 VSS.n1178 VSS.n1177 585
R511 VSS.n1179 VSS.n1178 585
R512 VSS.n1168 VSS.n1037 585
R513 VSS.n1037 VSS.n1036 585
R514 VSS.n1167 VSS.n1166 585
R515 VSS.n1166 VSS.n1165 585
R516 VSS.n1040 VSS.n1039 585
R517 VSS.n1041 VSS.n1040 585
R518 VSS.n1158 VSS.n1157 585
R519 VSS.n1159 VSS.n1158 585
R520 VSS.n1156 VSS.n1045 585
R521 VSS.n1050 VSS.n1045 585
R522 VSS.n1155 VSS.n1154 585
R523 VSS.n1154 VSS.n1153 585
R524 VSS.n1047 VSS.n1046 585
R525 VSS.n1048 VSS.n1047 585
R526 VSS.n1074 VSS.n1073 585
R527 VSS.n1076 VSS.n1075 585
R528 VSS.n1078 VSS.n1077 585
R529 VSS.n1080 VSS.n1079 585
R530 VSS.n1082 VSS.n1081 585
R531 VSS.n1084 VSS.n1083 585
R532 VSS.n1086 VSS.n1085 585
R533 VSS.n1088 VSS.n1087 585
R534 VSS.n1090 VSS.n1089 585
R535 VSS.n1092 VSS.n1091 585
R536 VSS.n1094 VSS.n1093 585
R537 VSS.n1096 VSS.n1095 585
R538 VSS.n1098 VSS.n1097 585
R539 VSS.n1100 VSS.n1099 585
R540 VSS.n1102 VSS.n1101 585
R541 VSS.n1104 VSS.n1103 585
R542 VSS.n1106 VSS.n1105 585
R543 VSS.n1108 VSS.n1107 585
R544 VSS.n1110 VSS.n1109 585
R545 VSS.n1112 VSS.n1111 585
R546 VSS.n1114 VSS.n1113 585
R547 VSS.n1116 VSS.n1115 585
R548 VSS.n1118 VSS.n1117 585
R549 VSS.n1120 VSS.n1119 585
R550 VSS.n1122 VSS.n1121 585
R551 VSS.n1124 VSS.n1123 585
R552 VSS.n1126 VSS.n1125 585
R553 VSS.n1128 VSS.n1127 585
R554 VSS.n1130 VSS.n1129 585
R555 VSS.n1132 VSS.n1131 585
R556 VSS.n1134 VSS.n1133 585
R557 VSS.n1136 VSS.n1135 585
R558 VSS.n1138 VSS.n1137 585
R559 VSS.n1140 VSS.n1139 585
R560 VSS.n1142 VSS.n1141 585
R561 VSS.n1143 VSS.n1072 585
R562 VSS.n1145 VSS.n1144 585
R563 VSS.n1053 VSS.n1052 585
R564 VSS.n1149 VSS.n1148 585
R565 VSS.n1148 VSS.n1147 585
R566 VSS.n1150 VSS.n1051 585
R567 VSS.n1051 VSS.n1048 585
R568 VSS.n1152 VSS.n1151 585
R569 VSS.n1153 VSS.n1152 585
R570 VSS.n1044 VSS.n1043 585
R571 VSS.n1050 VSS.n1044 585
R572 VSS.n1161 VSS.n1160 585
R573 VSS.n1160 VSS.n1159 585
R574 VSS.n1162 VSS.n1042 585
R575 VSS.n1042 VSS.n1041 585
R576 VSS.n1164 VSS.n1163 585
R577 VSS.n1165 VSS.n1164 585
R578 VSS.n1035 VSS.n1034 585
R579 VSS.n1036 VSS.n1035 585
R580 VSS.n1181 VSS.n1180 585
R581 VSS.n1180 VSS.n1179 585
R582 VSS.n1182 VSS.n1033 585
R583 VSS.n1033 VSS.n1031 585
R584 VSS.n1184 VSS.n1183 585
R585 VSS.n1185 VSS.n1184 585
R586 VSS.n1025 VSS.n1024 585
R587 VSS.n1026 VSS.n1025 585
R588 VSS.n1433 VSS.n1432 585
R589 VSS.n1432 VSS.n1431 585
R590 VSS.n1434 VSS.n1022 585
R591 VSS.n1022 VSS.n1019 585
R592 VSS.n1437 VSS.n1436 585
R593 VSS.n1438 VSS.n1437 585
R594 VSS.n1435 VSS.n1023 585
R595 VSS.n1023 VSS.n1013 585
R596 VSS.n1007 VSS.n1006 585
R597 VSS.n1447 VSS.n1007 585
R598 VSS.n1495 VSS.n1494 585
R599 VSS.n1494 VSS.n1493 585
R600 VSS.n1496 VSS.n1004 585
R601 VSS.n1491 VSS.n1004 585
R602 VSS.n1499 VSS.n1498 585
R603 VSS.n1500 VSS.n1499 585
R604 VSS.n1497 VSS.n1005 585
R605 VSS.n1005 VSS.n995 585
R606 VSS.n989 VSS.n988 585
R607 VSS.n996 VSS.n989 585
R608 VSS.n1519 VSS.n1518 585
R609 VSS.n1518 VSS.n1517 585
R610 VSS.n1520 VSS.n986 585
R611 VSS.n986 VSS.n982 585
R612 VSS.n1523 VSS.n1522 585
R613 VSS.n1524 VSS.n1523 585
R614 VSS.n1521 VSS.n987 585
R615 VSS.n987 VSS.n978 585
R616 VSS.n965 VSS.n964 585
R617 VSS.n1476 VSS.n965 585
R618 VSS.n1564 VSS.n1563 585
R619 VSS.n1563 VSS.n1562 585
R620 VSS.n1565 VSS.n963 585
R621 VSS.n969 VSS.n963 585
R622 VSS.n1567 VSS.n1566 585
R623 VSS.n1568 VSS.n1567 585
R624 VSS.n951 VSS.n950 585
R625 VSS.n974 VSS.n951 585
R626 VSS.n1644 VSS.n1643 585
R627 VSS.n1643 VSS.n1642 585
R628 VSS.n1645 VSS.n949 585
R629 VSS.n956 VSS.n949 585
R630 VSS.n1647 VSS.n1646 585
R631 VSS.n1648 VSS.n1647 585
R632 VSS.n930 VSS.n929 585
R633 VSS.n1657 VSS.n930 585
R634 VSS.n1668 VSS.n1667 585
R635 VSS.n1667 VSS.n1666 585
R636 VSS.n1669 VSS.n928 585
R637 VSS.n935 VSS.n928 585
R638 VSS.n1671 VSS.n1670 585
R639 VSS.n1672 VSS.n1671 585
R640 VSS.n909 VSS.n908 585
R641 VSS.n1681 VSS.n909 585
R642 VSS.n1692 VSS.n1691 585
R643 VSS.n1691 VSS.n1690 585
R644 VSS.n1693 VSS.n906 585
R645 VSS.n906 VSS.n903 585
R646 VSS.n1696 VSS.n1695 585
R647 VSS.n1697 VSS.n1696 585
R648 VSS.n1694 VSS.n907 585
R649 VSS.n907 VSS.n735 585
R650 VSS.n794 VSS.n792 585
R651 VSS.n898 VSS.n792 585
R652 VSS.n2044 VSS.n2043 585
R653 VSS.n2045 VSS.n2044 585
R654 VSS.n2042 VSS.n793 585
R655 VSS.n1788 VSS.n793 585
R656 VSS.n2041 VSS.n2040 585
R657 VSS.n2040 VSS.n2039 585
R658 VSS.n796 VSS.n795 585
R659 VSS.n800 VSS.n796 585
R660 VSS.n822 VSS.n821 585
R661 VSS.n822 VSS.n806 585
R662 VSS.n824 VSS.n823 585
R663 VSS.n823 VSS.n809 585
R664 VSS.n825 VSS.n819 585
R665 VSS.n1799 VSS.n819 585
R666 VSS.n2023 VSS.n2022 585
R667 VSS.n2024 VSS.n2023 585
R668 VSS.n2021 VSS.n820 585
R669 VSS.n1992 VSS.n820 585
R670 VSS.n2020 VSS.n2019 585
R671 VSS.n2019 VSS.n2018 585
R672 VSS.n831 VSS.n826 585
R673 VSS.n2012 VSS.n831 585
R674 VSS.n830 VSS.n829 585
R675 VSS.n830 VSS.n332 585
R676 VSS.n828 VSS.n827 585
R677 VSS.n827 VSS.n334 585
R678 VSS.n346 VSS.n344 585
R679 VSS.n2002 VSS.n344 585
R680 VSS.n2304 VSS.n2303 585
R681 VSS.n2305 VSS.n2304 585
R682 VSS.n2302 VSS.n345 585
R683 VSS.n2250 VSS.n345 585
R684 VSS.n2301 VSS.n2300 585
R685 VSS.n2300 VSS.n2299 585
R686 VSS.n348 VSS.n347 585
R687 VSS.n360 VSS.n348 585
R688 VSS.n2150 VSS.n2149 585
R689 VSS.n2151 VSS.n2150 585
R690 VSS.n2050 VSS.n737 585
R691 VSS.n2049 VSS.n2048 585
R692 VSS.n740 VSS.n739 585
R693 VSS.n2046 VSS.n740 585
R694 VSS.n753 VSS.n752 585
R695 VSS.n755 VSS.n754 585
R696 VSS.n757 VSS.n756 585
R697 VSS.n759 VSS.n758 585
R698 VSS.n761 VSS.n760 585
R699 VSS.n763 VSS.n762 585
R700 VSS.n765 VSS.n764 585
R701 VSS.n767 VSS.n766 585
R702 VSS.n769 VSS.n768 585
R703 VSS.n771 VSS.n770 585
R704 VSS.n773 VSS.n772 585
R705 VSS.n775 VSS.n774 585
R706 VSS.n777 VSS.n776 585
R707 VSS.n779 VSS.n778 585
R708 VSS.n781 VSS.n780 585
R709 VSS.n783 VSS.n782 585
R710 VSS.n785 VSS.n784 585
R711 VSS.n786 VSS.n751 585
R712 VSS.n788 VSS.n787 585
R713 VSS.n733 VSS.n731 585
R714 VSS.n2055 VSS.n2054 585
R715 VSS.n2054 VSS.n2053 585
R716 VSS.n732 VSS.n730 585
R717 VSS.n1698 VSS.n732 585
R718 VSS.n914 VSS.n913 585
R719 VSS.n1688 VSS.n914 585
R720 VSS.n1581 VSS.n1580 585
R721 VSS.n1580 VSS.n910 585
R722 VSS.n1582 VSS.n919 585
R723 VSS.n1682 VSS.n919 585
R724 VSS.n1583 VSS.n926 585
R725 VSS.n1673 VSS.n926 585
R726 VSS.n1584 VSS.n934 585
R727 VSS.n1664 VSS.n934 585
R728 VSS.n1586 VSS.n1585 585
R729 VSS.n1585 VSS.n931 585
R730 VSS.n1587 VSS.n940 585
R731 VSS.n1658 VSS.n940 585
R732 VSS.n1588 VSS.n947 585
R733 VSS.n1649 VSS.n947 585
R734 VSS.n1589 VSS.n955 585
R735 VSS.n1640 VSS.n955 585
R736 VSS.n1591 VSS.n1590 585
R737 VSS.n1591 VSS.n952 585
R738 VSS.n1593 VSS.n1592 585
R739 VSS.n1595 VSS.n1594 585
R740 VSS.n1597 VSS.n1596 585
R741 VSS.n1599 VSS.n1598 585
R742 VSS.n1601 VSS.n1600 585
R743 VSS.n1603 VSS.n1602 585
R744 VSS.n1605 VSS.n1604 585
R745 VSS.n1607 VSS.n1606 585
R746 VSS.n1609 VSS.n1608 585
R747 VSS.n1611 VSS.n1610 585
R748 VSS.n1613 VSS.n1612 585
R749 VSS.n1615 VSS.n1614 585
R750 VSS.n1617 VSS.n1616 585
R751 VSS.n1619 VSS.n1618 585
R752 VSS.n1621 VSS.n1620 585
R753 VSS.n1623 VSS.n1622 585
R754 VSS.n1625 VSS.n1624 585
R755 VSS.n1627 VSS.n1626 585
R756 VSS.n1629 VSS.n1628 585
R757 VSS.n1630 VSS.n1579 585
R758 VSS.n1632 VSS.n1631 585
R759 VSS.n959 VSS.n958 585
R760 VSS.n1636 VSS.n1635 585
R761 VSS.n1635 VSS.n1634 585
R762 VSS.n1637 VSS.n957 585
R763 VSS.n957 VSS.n952 585
R764 VSS.n1639 VSS.n1638 585
R765 VSS.n1640 VSS.n1639 585
R766 VSS.n938 VSS.n937 585
R767 VSS.n1649 VSS.n938 585
R768 VSS.n1660 VSS.n1659 585
R769 VSS.n1659 VSS.n1658 585
R770 VSS.n1661 VSS.n936 585
R771 VSS.n936 VSS.n931 585
R772 VSS.n1663 VSS.n1662 585
R773 VSS.n1664 VSS.n1663 585
R774 VSS.n917 VSS.n916 585
R775 VSS.n1673 VSS.n917 585
R776 VSS.n1684 VSS.n1683 585
R777 VSS.n1683 VSS.n1682 585
R778 VSS.n1685 VSS.n915 585
R779 VSS.n915 VSS.n910 585
R780 VSS.n1687 VSS.n1686 585
R781 VSS.n1688 VSS.n1687 585
R782 VSS.n738 VSS.n736 585
R783 VSS.n1698 VSS.n736 585
R784 VSS.n2052 VSS.n2051 585
R785 VSS.n2053 VSS.n2052 585
R786 VSS.n2296 VSS.n2295 585
R787 VSS.n2294 VSS.n362 585
R788 VSS.n2293 VSS.n361 585
R789 VSS.n2298 VSS.n361 585
R790 VSS.n2292 VSS.n2291 585
R791 VSS.n2290 VSS.n2289 585
R792 VSS.n2288 VSS.n2287 585
R793 VSS.n2286 VSS.n2285 585
R794 VSS.n2284 VSS.n2283 585
R795 VSS.n2282 VSS.n2281 585
R796 VSS.n2280 VSS.n2279 585
R797 VSS.n2278 VSS.n2277 585
R798 VSS.n2276 VSS.n2275 585
R799 VSS.n2274 VSS.n2273 585
R800 VSS.n2272 VSS.n2271 585
R801 VSS.n2270 VSS.n2269 585
R802 VSS.n2268 VSS.n2267 585
R803 VSS.n2266 VSS.n2265 585
R804 VSS.n2264 VSS.n2263 585
R805 VSS.n2262 VSS.n2261 585
R806 VSS.n2260 VSS.n2259 585
R807 VSS.n2258 VSS.n2257 585
R808 VSS.n2256 VSS.n2255 585
R809 VSS.n2254 VSS.n2253 585
R810 VSS.n2252 VSS.n363 585
R811 VSS.n2252 VSS.n2251 585
R812 VSS.n837 VSS.n341 585
R813 VSS.n2306 VSS.n341 585
R814 VSS.n2005 VSS.n2004 585
R815 VSS.n2004 VSS.n2003 585
R816 VSS.n2007 VSS.n333 585
R817 VSS.n2312 VSS.n333 585
R818 VSS.n2010 VSS.n2009 585
R819 VSS.n2011 VSS.n2010 585
R820 VSS.n836 VSS.n834 585
R821 VSS.n2017 VSS.n834 585
R822 VSS.n1772 VSS.n1771 585
R823 VSS.n1772 VSS.n832 585
R824 VSS.n1774 VSS.n1773 585
R825 VSS.n1773 VSS.n818 585
R826 VSS.n1775 VSS.n816 585
R827 VSS.n2025 VSS.n816 585
R828 VSS.n1776 VSS.n892 585
R829 VSS.n1800 VSS.n892 585
R830 VSS.n1777 VSS.n808 585
R831 VSS.n2031 VSS.n808 585
R832 VSS.n1779 VSS.n1778 585
R833 VSS.n1780 VSS.n1779 585
R834 VSS.n1770 VSS.n1714 585
R835 VSS.n1769 VSS.n1768 585
R836 VSS.n1766 VSS.n1715 585
R837 VSS.n1764 VSS.n1763 585
R838 VSS.n1762 VSS.n1716 585
R839 VSS.n1761 VSS.n1760 585
R840 VSS.n1758 VSS.n1717 585
R841 VSS.n1756 VSS.n1755 585
R842 VSS.n1754 VSS.n1718 585
R843 VSS.n1753 VSS.n1752 585
R844 VSS.n1750 VSS.n1719 585
R845 VSS.n1748 VSS.n1747 585
R846 VSS.n1746 VSS.n1720 585
R847 VSS.n1745 VSS.n1744 585
R848 VSS.n1742 VSS.n1721 585
R849 VSS.n1740 VSS.n1739 585
R850 VSS.n1738 VSS.n1722 585
R851 VSS.n1737 VSS.n1736 585
R852 VSS.n1734 VSS.n1723 585
R853 VSS.n1732 VSS.n1731 585
R854 VSS.n1730 VSS.n1724 585
R855 VSS.n1729 VSS.n1728 585
R856 VSS.n1726 VSS.n1725 585
R857 VSS.n1726 VSS.n797 585
R858 VSS.n812 VSS.n810 585
R859 VSS.n1780 VSS.n810 585
R860 VSS.n2030 VSS.n2029 585
R861 VSS.n2031 VSS.n2030 585
R862 VSS.n2028 VSS.n811 585
R863 VSS.n1800 VSS.n811 585
R864 VSS.n2027 VSS.n2026 585
R865 VSS.n2026 VSS.n2025 585
R866 VSS.n814 VSS.n813 585
R867 VSS.n818 VSS.n814 585
R868 VSS.n2014 VSS.n2013 585
R869 VSS.n2013 VSS.n832 585
R870 VSS.n2016 VSS.n2015 585
R871 VSS.n2017 VSS.n2016 585
R872 VSS.n337 VSS.n335 585
R873 VSS.n2011 VSS.n335 585
R874 VSS.n2311 VSS.n2310 585
R875 VSS.n2312 VSS.n2311 585
R876 VSS.n2309 VSS.n336 585
R877 VSS.n2003 VSS.n336 585
R878 VSS.n2308 VSS.n2307 585
R879 VSS.n2307 VSS.n2306 585
R880 VSS.n339 VSS.n338 585
R881 VSS.n2251 VSS.n339 585
R882 VSS.n2117 VSS.n2116 585
R883 VSS.n2115 VSS.n596 585
R884 VSS.n2114 VSS.n595 585
R885 VSS.n2119 VSS.n595 585
R886 VSS.n2113 VSS.n2112 585
R887 VSS.n2111 VSS.n2110 585
R888 VSS.n2109 VSS.n2108 585
R889 VSS.n2107 VSS.n2106 585
R890 VSS.n2105 VSS.n2104 585
R891 VSS.n2103 VSS.n2102 585
R892 VSS.n2101 VSS.n2100 585
R893 VSS.n2099 VSS.n2098 585
R894 VSS.n2097 VSS.n2096 585
R895 VSS.n2095 VSS.n2094 585
R896 VSS.n2093 VSS.n2092 585
R897 VSS.n2091 VSS.n2090 585
R898 VSS.n2089 VSS.n2088 585
R899 VSS.n2087 VSS.n2086 585
R900 VSS.n2085 VSS.n2084 585
R901 VSS.n2083 VSS.n2082 585
R902 VSS.n2081 VSS.n2080 585
R903 VSS.n2079 VSS.n2078 585
R904 VSS.n2077 VSS.n2076 585
R905 VSS.n2075 VSS.n2074 585
R906 VSS.n2073 VSS.n584 585
R907 VSS.n2120 VSS.n584 585
R908 VSS.n2072 VSS.n583 585
R909 VSS.n2121 VSS.n583 585
R910 VSS.n2071 VSS.n2070 585
R911 VSS.n2070 VSS.n579 585
R912 VSS.n2069 VSS.n578 585
R913 VSS.n2127 VSS.n578 585
R914 VSS.n2068 VSS.n577 585
R915 VSS.n2128 VSS.n577 585
R916 VSS.n2067 VSS.n576 585
R917 VSS.n2129 VSS.n576 585
R918 VSS.n2066 VSS.n2065 585
R919 VSS.n2065 VSS.n572 585
R920 VSS.n2064 VSS.n571 585
R921 VSS.n2135 VSS.n571 585
R922 VSS.n2063 VSS.n570 585
R923 VSS.n2136 VSS.n570 585
R924 VSS.n2062 VSS.n569 585
R925 VSS.n2137 VSS.n569 585
R926 VSS.n598 VSS.n597 585
R927 VSS.n597 VSS.n563 585
R928 VSS.n654 VSS.n562 585
R929 VSS.n2143 VSS.n562 585
R930 VSS.n653 VSS.n652 585
R931 VSS.n650 VSS.n599 585
R932 VSS.n649 VSS.n648 585
R933 VSS.n647 VSS.n646 585
R934 VSS.n645 VSS.n601 585
R935 VSS.n643 VSS.n642 585
R936 VSS.n641 VSS.n602 585
R937 VSS.n640 VSS.n639 585
R938 VSS.n637 VSS.n603 585
R939 VSS.n635 VSS.n634 585
R940 VSS.n633 VSS.n604 585
R941 VSS.n632 VSS.n631 585
R942 VSS.n629 VSS.n605 585
R943 VSS.n627 VSS.n626 585
R944 VSS.n625 VSS.n606 585
R945 VSS.n624 VSS.n623 585
R946 VSS.n621 VSS.n607 585
R947 VSS.n619 VSS.n618 585
R948 VSS.n617 VSS.n608 585
R949 VSS.n616 VSS.n615 585
R950 VSS.n613 VSS.n609 585
R951 VSS.n611 VSS.n610 585
R952 VSS.n566 VSS.n564 585
R953 VSS.n564 VSS.n367 585
R954 VSS.n2142 VSS.n2141 585
R955 VSS.n2143 VSS.n2142 585
R956 VSS.n2140 VSS.n565 585
R957 VSS.n565 VSS.n563 585
R958 VSS.n2139 VSS.n2138 585
R959 VSS.n2138 VSS.n2137 585
R960 VSS.n568 VSS.n567 585
R961 VSS.n2136 VSS.n568 585
R962 VSS.n2134 VSS.n2133 585
R963 VSS.n2135 VSS.n2134 585
R964 VSS.n2132 VSS.n573 585
R965 VSS.n573 VSS.n572 585
R966 VSS.n2131 VSS.n2130 585
R967 VSS.n2130 VSS.n2129 585
R968 VSS.n575 VSS.n574 585
R969 VSS.n2128 VSS.n575 585
R970 VSS.n2126 VSS.n2125 585
R971 VSS.n2127 VSS.n2126 585
R972 VSS.n2124 VSS.n580 585
R973 VSS.n580 VSS.n579 585
R974 VSS.n2123 VSS.n2122 585
R975 VSS.n2122 VSS.n2121 585
R976 VSS.n582 VSS.n581 585
R977 VSS.n2120 VSS.n582 585
R978 VSS.n2248 VSS.n2247 585
R979 VSS.n2249 VSS.n2248 585
R980 VSS.n2163 VSS.n2158 585
R981 VSS.n2158 VSS.n343 585
R982 VSS.n2162 VSS.n2161 585
R983 VSS.n2161 VSS.n340 585
R984 VSS.n2160 VSS.n331 585
R985 VSS.n838 VSS.n331 585
R986 VSS.n2314 VSS.n329 585
R987 VSS.n2314 VSS.n2313 585
R988 VSS.n1418 VSS.n1028 585
R989 VSS.n1417 VSS.n1416 585
R990 VSS.n1030 VSS.n1029 585
R991 VSS.n1412 VSS.n1411 585
R992 VSS.n1410 VSS.n1231 585
R993 VSS.n1409 VSS.n1408 585
R994 VSS.n1407 VSS.n1406 585
R995 VSS.n1405 VSS.n1404 585
R996 VSS.n1403 VSS.n1402 585
R997 VSS.n1401 VSS.n1400 585
R998 VSS.n1399 VSS.n1398 585
R999 VSS.n1397 VSS.n1396 585
R1000 VSS.n1395 VSS.n1394 585
R1001 VSS.n1393 VSS.n1392 585
R1002 VSS.n1391 VSS.n1390 585
R1003 VSS.n1389 VSS.n1388 585
R1004 VSS.n1387 VSS.n1386 585
R1005 VSS.n1385 VSS.n1384 585
R1006 VSS.n1383 VSS.n1382 585
R1007 VSS.n1381 VSS.n1380 585
R1008 VSS.n1379 VSS.n1378 585
R1009 VSS.n1377 VSS.n1376 585
R1010 VSS.n1375 VSS.n1374 585
R1011 VSS.n1373 VSS.n1372 585
R1012 VSS.n1371 VSS.n1370 585
R1013 VSS.n1369 VSS.n1368 585
R1014 VSS.n1367 VSS.n1366 585
R1015 VSS.n1365 VSS.n1364 585
R1016 VSS.n1363 VSS.n1362 585
R1017 VSS.n1361 VSS.n1360 585
R1018 VSS.n1359 VSS.n1358 585
R1019 VSS.n1357 VSS.n1356 585
R1020 VSS.n1355 VSS.n1354 585
R1021 VSS.n1353 VSS.n1352 585
R1022 VSS.n1351 VSS.n1350 585
R1023 VSS.n1349 VSS.n1348 585
R1024 VSS.n1347 VSS.n1346 585
R1025 VSS.n1345 VSS.n1344 585
R1026 VSS.n1343 VSS.n1342 585
R1027 VSS.n1341 VSS.n1340 585
R1028 VSS.n1339 VSS.n1338 585
R1029 VSS.n1337 VSS.n1336 585
R1030 VSS.n1335 VSS.n1334 585
R1031 VSS.n1333 VSS.n1332 585
R1032 VSS.n1331 VSS.n1330 585
R1033 VSS.n1329 VSS.n1328 585
R1034 VSS.n1327 VSS.n1326 585
R1035 VSS.n1325 VSS.n1324 585
R1036 VSS.n1323 VSS.n1322 585
R1037 VSS.n1321 VSS.n1320 585
R1038 VSS.n1319 VSS.n1318 585
R1039 VSS.n1317 VSS.n1316 585
R1040 VSS.n1315 VSS.n1314 585
R1041 VSS.n1313 VSS.n1312 585
R1042 VSS.n1311 VSS.n1310 585
R1043 VSS.n1309 VSS.n1308 585
R1044 VSS.n1307 VSS.n1306 585
R1045 VSS.n1305 VSS.n1304 585
R1046 VSS.n1303 VSS.n1302 585
R1047 VSS.n1301 VSS.n1300 585
R1048 VSS.n1299 VSS.n1298 585
R1049 VSS.n1297 VSS.n1296 585
R1050 VSS.n1295 VSS.n1294 585
R1051 VSS.n1293 VSS.n1292 585
R1052 VSS.n1291 VSS.n1290 585
R1053 VSS.n1289 VSS.n1288 585
R1054 VSS.n1287 VSS.n1286 585
R1055 VSS.n1285 VSS.n1284 585
R1056 VSS.n1283 VSS.n1282 585
R1057 VSS.n1281 VSS.n1280 585
R1058 VSS.n1279 VSS.n1278 585
R1059 VSS.n1277 VSS.n1276 585
R1060 VSS.n1275 VSS.n1274 585
R1061 VSS.n1273 VSS.n1272 585
R1062 VSS.n1271 VSS.n1270 585
R1063 VSS.n1269 VSS.n1268 585
R1064 VSS.n1267 VSS.n1266 585
R1065 VSS.n1265 VSS.n1264 585
R1066 VSS.n1263 VSS.n1262 585
R1067 VSS.n1261 VSS.n1260 585
R1068 VSS.n1259 VSS.n1258 585
R1069 VSS.n1257 VSS.n1256 585
R1070 VSS.n1255 VSS.n1254 585
R1071 VSS.n1253 VSS.n1252 585
R1072 VSS.n1251 VSS.n1250 585
R1073 VSS.n1249 VSS.n1248 585
R1074 VSS.n1247 VSS.n1246 585
R1075 VSS.n1245 VSS.n1244 585
R1076 VSS.n1243 VSS.n1242 585
R1077 VSS.n1241 VSS.n1240 585
R1078 VSS.n1239 VSS.n1238 585
R1079 VSS.n1237 VSS.n1236 585
R1080 VSS.n1235 VSS.n1234 585
R1081 VSS.n1233 VSS.n1232 585
R1082 VSS.n1018 VSS.n1017 585
R1083 VSS.n1430 VSS.n1018 585
R1084 VSS.n1441 VSS.n1440 585
R1085 VSS.n1440 VSS.n1439 585
R1086 VSS.n1442 VSS.n1015 585
R1087 VSS.n1424 VSS.n1015 585
R1088 VSS.n1445 VSS.n1444 585
R1089 VSS.n1446 VSS.n1445 585
R1090 VSS.n1443 VSS.n1016 585
R1091 VSS.n1016 VSS.n1008 585
R1092 VSS.n1000 VSS.n999 585
R1093 VSS.n1492 VSS.n1000 585
R1094 VSS.n1503 VSS.n1502 585
R1095 VSS.n1502 VSS.n1501 585
R1096 VSS.n1504 VSS.n997 585
R1097 VSS.n1003 VSS.n997 585
R1098 VSS.n1507 VSS.n1506 585
R1099 VSS.n1508 VSS.n1507 585
R1100 VSS.n1505 VSS.n998 585
R1101 VSS.n998 VSS.n990 585
R1102 VSS.n981 VSS.n980 585
R1103 VSS.n1516 VSS.n981 585
R1104 VSS.n1527 VSS.n1526 585
R1105 VSS.n1526 VSS.n1525 585
R1106 VSS.n1528 VSS.n979 585
R1107 VSS.n985 VSS.n979 585
R1108 VSS.n1530 VSS.n1529 585
R1109 VSS.n1531 VSS.n1530 585
R1110 VSS.n972 VSS.n970 585
R1111 VSS.n970 VSS.n966 585
R1112 VSS.n1560 VSS.n1559 585
R1113 VSS.n1561 VSS.n1560 585
R1114 VSS.n1558 VSS.n971 585
R1115 VSS.n971 VSS.n960 585
R1116 VSS.n1557 VSS.n1556 585
R1117 VSS.n1556 VSS.n962 585
R1118 VSS.n1555 VSS.n973 585
R1119 VSS.n1555 VSS.n1554 585
R1120 VSS.n945 VSS.n944 585
R1121 VSS.n1641 VSS.n945 585
R1122 VSS.n1652 VSS.n1651 585
R1123 VSS.n1651 VSS.n1650 585
R1124 VSS.n1653 VSS.n943 585
R1125 VSS.n943 VSS.n939 585
R1126 VSS.n1655 VSS.n1654 585
R1127 VSS.n1656 VSS.n1655 585
R1128 VSS.n924 VSS.n923 585
R1129 VSS.n1665 VSS.n924 585
R1130 VSS.n1676 VSS.n1675 585
R1131 VSS.n1675 VSS.n1674 585
R1132 VSS.n1677 VSS.n922 585
R1133 VSS.n922 VSS.n918 585
R1134 VSS.n1679 VSS.n1678 585
R1135 VSS.n1680 VSS.n1679 585
R1136 VSS.n902 VSS.n901 585
R1137 VSS.n1689 VSS.n902 585
R1138 VSS.n1701 VSS.n1700 585
R1139 VSS.n1700 VSS.n1699 585
R1140 VSS.n1702 VSS.n899 585
R1141 VSS.n899 VSS.n734 585
R1142 VSS.n1707 VSS.n1706 585
R1143 VSS.n1708 VSS.n1707 585
R1144 VSS.n1705 VSS.n900 585
R1145 VSS.n900 VSS.n741 585
R1146 VSS.n1704 VSS.n1703 585
R1147 VSS.n1703 VSS.n791 585
R1148 VSS.n803 VSS.n801 585
R1149 VSS.n1787 VSS.n801 585
R1150 VSS.n2037 VSS.n2036 585
R1151 VSS.n2038 VSS.n2037 585
R1152 VSS.n2035 VSS.n802 585
R1153 VSS.n1781 VSS.n802 585
R1154 VSS.n2034 VSS.n2033 585
R1155 VSS.n2033 VSS.n2032 585
R1156 VSS.n805 VSS.n804 585
R1157 VSS.n1801 VSS.n805 585
R1158 VSS.n890 VSS.n889 585
R1159 VSS.n889 VSS.n815 585
R1160 VSS.n1989 VSS.n1988 585
R1161 VSS.n1987 VSS.n888 585
R1162 VSS.n1986 VSS.n887 585
R1163 VSS.n1991 VSS.n887 585
R1164 VSS.n1985 VSS.n1984 585
R1165 VSS.n1983 VSS.n1982 585
R1166 VSS.n1981 VSS.n1980 585
R1167 VSS.n1979 VSS.n1978 585
R1168 VSS.n1977 VSS.n1976 585
R1169 VSS.n1975 VSS.n1974 585
R1170 VSS.n1973 VSS.n1972 585
R1171 VSS.n1971 VSS.n1970 585
R1172 VSS.n1969 VSS.n1968 585
R1173 VSS.n1967 VSS.n1966 585
R1174 VSS.n1965 VSS.n1964 585
R1175 VSS.n1963 VSS.n1962 585
R1176 VSS.n1961 VSS.n1960 585
R1177 VSS.n1959 VSS.n1958 585
R1178 VSS.n1957 VSS.n1956 585
R1179 VSS.n1955 VSS.n1954 585
R1180 VSS.n1953 VSS.n1952 585
R1181 VSS.n1951 VSS.n1950 585
R1182 VSS.n1949 VSS.n1948 585
R1183 VSS.n1947 VSS.n1946 585
R1184 VSS.n1945 VSS.n1944 585
R1185 VSS.n1943 VSS.n1942 585
R1186 VSS.n1941 VSS.n1940 585
R1187 VSS.n1939 VSS.n1938 585
R1188 VSS.n1937 VSS.n1936 585
R1189 VSS.n1935 VSS.n1934 585
R1190 VSS.n1933 VSS.n1932 585
R1191 VSS.n1931 VSS.n1930 585
R1192 VSS.n1929 VSS.n1928 585
R1193 VSS.n1927 VSS.n1926 585
R1194 VSS.n1925 VSS.n1924 585
R1195 VSS.n1923 VSS.n1922 585
R1196 VSS.n1921 VSS.n1920 585
R1197 VSS.n1919 VSS.n1918 585
R1198 VSS.n1917 VSS.n1916 585
R1199 VSS.n1915 VSS.n1914 585
R1200 VSS.n1913 VSS.n1912 585
R1201 VSS.n1911 VSS.n1910 585
R1202 VSS.n1909 VSS.n1908 585
R1203 VSS.n1907 VSS.n1906 585
R1204 VSS.n1905 VSS.n1904 585
R1205 VSS.n1903 VSS.n1902 585
R1206 VSS.n1901 VSS.n1900 585
R1207 VSS.n1899 VSS.n1898 585
R1208 VSS.n1897 VSS.n1896 585
R1209 VSS.n1895 VSS.n1894 585
R1210 VSS.n1893 VSS.n1892 585
R1211 VSS.n1891 VSS.n1890 585
R1212 VSS.n1889 VSS.n1888 585
R1213 VSS.n1887 VSS.n1886 585
R1214 VSS.n1885 VSS.n1884 585
R1215 VSS.n1883 VSS.n1882 585
R1216 VSS.n1881 VSS.n1880 585
R1217 VSS.n1879 VSS.n1878 585
R1218 VSS.n1877 VSS.n1876 585
R1219 VSS.n1875 VSS.n1874 585
R1220 VSS.n1873 VSS.n1872 585
R1221 VSS.n1871 VSS.n1870 585
R1222 VSS.n1869 VSS.n1868 585
R1223 VSS.n1867 VSS.n1866 585
R1224 VSS.n1865 VSS.n1864 585
R1225 VSS.n1863 VSS.n1862 585
R1226 VSS.n1861 VSS.n1860 585
R1227 VSS.n1859 VSS.n1858 585
R1228 VSS.n1857 VSS.n1856 585
R1229 VSS.n1855 VSS.n1854 585
R1230 VSS.n1853 VSS.n1852 585
R1231 VSS.n1851 VSS.n1850 585
R1232 VSS.n1849 VSS.n1848 585
R1233 VSS.n1847 VSS.n1846 585
R1234 VSS.n1845 VSS.n1844 585
R1235 VSS.n1843 VSS.n1842 585
R1236 VSS.n1841 VSS.n1840 585
R1237 VSS.n1839 VSS.n1838 585
R1238 VSS.n1837 VSS.n1836 585
R1239 VSS.n1835 VSS.n1834 585
R1240 VSS.n1833 VSS.n1832 585
R1241 VSS.n1831 VSS.n1830 585
R1242 VSS.n1829 VSS.n1828 585
R1243 VSS.n1827 VSS.n1826 585
R1244 VSS.n1825 VSS.n1824 585
R1245 VSS.n1823 VSS.n1822 585
R1246 VSS.n1821 VSS.n1820 585
R1247 VSS.n1819 VSS.n1818 585
R1248 VSS.n1817 VSS.n1816 585
R1249 VSS.n1815 VSS.n1814 585
R1250 VSS.n1813 VSS.n1812 585
R1251 VSS.n1811 VSS.n1810 585
R1252 VSS.n1809 VSS.n1808 585
R1253 VSS.n1807 VSS.n1806 585
R1254 VSS.n1805 VSS.n886 585
R1255 VSS.n1991 VSS.n886 585
R1256 VSS.n1804 VSS.n1803 585
R1257 VSS.n1803 VSS.n815 585
R1258 VSS.n1802 VSS.n891 585
R1259 VSS.n1802 VSS.n1801 585
R1260 VSS.n1713 VSS.n807 585
R1261 VSS.n2032 VSS.n807 585
R1262 VSS.n1783 VSS.n1782 585
R1263 VSS.n1782 VSS.n1781 585
R1264 VSS.n1784 VSS.n799 585
R1265 VSS.n2038 VSS.n799 585
R1266 VSS.n1786 VSS.n1785 585
R1267 VSS.n1787 VSS.n1786 585
R1268 VSS.n1712 VSS.n895 585
R1269 VSS.n895 VSS.n791 585
R1270 VSS.n1711 VSS.n1710 585
R1271 VSS.n1710 VSS.n741 585
R1272 VSS.n1709 VSS.n896 585
R1273 VSS.n1709 VSS.n1708 585
R1274 VSS.n1539 VSS.n897 585
R1275 VSS.n897 VSS.n734 585
R1276 VSS.n1540 VSS.n904 585
R1277 VSS.n1699 VSS.n904 585
R1278 VSS.n1541 VSS.n912 585
R1279 VSS.n1689 VSS.n912 585
R1280 VSS.n1542 VSS.n921 585
R1281 VSS.n1680 VSS.n921 585
R1282 VSS.n1544 VSS.n1543 585
R1283 VSS.n1543 VSS.n918 585
R1284 VSS.n1545 VSS.n925 585
R1285 VSS.n1674 VSS.n925 585
R1286 VSS.n1546 VSS.n933 585
R1287 VSS.n1665 VSS.n933 585
R1288 VSS.n1547 VSS.n942 585
R1289 VSS.n1656 VSS.n942 585
R1290 VSS.n1549 VSS.n1548 585
R1291 VSS.n1548 VSS.n939 585
R1292 VSS.n1550 VSS.n946 585
R1293 VSS.n1650 VSS.n946 585
R1294 VSS.n1551 VSS.n954 585
R1295 VSS.n1641 VSS.n954 585
R1296 VSS.n1553 VSS.n1552 585
R1297 VSS.n1554 VSS.n1553 585
R1298 VSS.n1538 VSS.n975 585
R1299 VSS.n975 VSS.n962 585
R1300 VSS.n1537 VSS.n1536 585
R1301 VSS.n1536 VSS.n960 585
R1302 VSS.n1535 VSS.n968 585
R1303 VSS.n1561 VSS.n968 585
R1304 VSS.n1534 VSS.n1533 585
R1305 VSS.n1533 VSS.n966 585
R1306 VSS.n1532 VSS.n976 585
R1307 VSS.n1532 VSS.n1531 585
R1308 VSS.n1512 VSS.n977 585
R1309 VSS.n985 VSS.n977 585
R1310 VSS.n1513 VSS.n983 585
R1311 VSS.n1525 VSS.n983 585
R1312 VSS.n1515 VSS.n1514 585
R1313 VSS.n1516 VSS.n1515 585
R1314 VSS.n1511 VSS.n992 585
R1315 VSS.n992 VSS.n990 585
R1316 VSS.n1510 VSS.n1509 585
R1317 VSS.n1509 VSS.n1508 585
R1318 VSS.n994 VSS.n993 585
R1319 VSS.n1003 VSS.n994 585
R1320 VSS.n1419 VSS.n1001 585
R1321 VSS.n1501 VSS.n1001 585
R1322 VSS.n1420 VSS.n1010 585
R1323 VSS.n1492 VSS.n1010 585
R1324 VSS.n1422 VSS.n1421 585
R1325 VSS.n1421 VSS.n1008 585
R1326 VSS.n1423 VSS.n1014 585
R1327 VSS.n1446 VSS.n1014 585
R1328 VSS.n1426 VSS.n1425 585
R1329 VSS.n1425 VSS.n1424 585
R1330 VSS.n1427 VSS.n1020 585
R1331 VSS.n1439 VSS.n1020 585
R1332 VSS.n1429 VSS.n1428 585
R1333 VSS.n1430 VSS.n1429 585
R1334 VSS.t123 VSS.n309 533.207
R1335 VSS.n2242 VSS.n2166 445.738
R1336 VSS.n2142 VSS.n565 394
R1337 VSS.n2138 VSS.n565 394
R1338 VSS.n2138 VSS.n568 394
R1339 VSS.n2134 VSS.n568 394
R1340 VSS.n2134 VSS.n573 394
R1341 VSS.n2130 VSS.n573 394
R1342 VSS.n2130 VSS.n575 394
R1343 VSS.n2126 VSS.n575 394
R1344 VSS.n2126 VSS.n580 394
R1345 VSS.n2122 VSS.n580 394
R1346 VSS.n2122 VSS.n582 394
R1347 VSS.n611 VSS.n564 394
R1348 VSS.n615 VSS.n613 394
R1349 VSS.n619 VSS.n608 394
R1350 VSS.n623 VSS.n621 394
R1351 VSS.n627 VSS.n606 394
R1352 VSS.n631 VSS.n629 394
R1353 VSS.n635 VSS.n604 394
R1354 VSS.n639 VSS.n637 394
R1355 VSS.n643 VSS.n602 394
R1356 VSS.n646 VSS.n645 394
R1357 VSS.n650 VSS.n649 394
R1358 VSS.n597 VSS.n562 394
R1359 VSS.n597 VSS.n569 394
R1360 VSS.n570 VSS.n569 394
R1361 VSS.n571 VSS.n570 394
R1362 VSS.n2065 VSS.n571 394
R1363 VSS.n2065 VSS.n576 394
R1364 VSS.n577 VSS.n576 394
R1365 VSS.n578 VSS.n577 394
R1366 VSS.n2070 VSS.n578 394
R1367 VSS.n2070 VSS.n583 394
R1368 VSS.n584 VSS.n583 394
R1369 VSS.n596 VSS.n595 394
R1370 VSS.n2112 VSS.n595 394
R1371 VSS.n2110 VSS.n2109 394
R1372 VSS.n2106 VSS.n2105 394
R1373 VSS.n2102 VSS.n2101 394
R1374 VSS.n2098 VSS.n2097 394
R1375 VSS.n2094 VSS.n2093 394
R1376 VSS.n2090 VSS.n2089 394
R1377 VSS.n2086 VSS.n2085 394
R1378 VSS.n2082 VSS.n2081 394
R1379 VSS.n2078 VSS.n2077 394
R1380 VSS.n2030 VSS.n810 394
R1381 VSS.n2030 VSS.n811 394
R1382 VSS.n2026 VSS.n811 394
R1383 VSS.n2026 VSS.n814 394
R1384 VSS.n2013 VSS.n814 394
R1385 VSS.n2016 VSS.n2013 394
R1386 VSS.n2016 VSS.n335 394
R1387 VSS.n2311 VSS.n335 394
R1388 VSS.n2311 VSS.n336 394
R1389 VSS.n2307 VSS.n336 394
R1390 VSS.n2307 VSS.n339 394
R1391 VSS.n1728 VSS.n1726 394
R1392 VSS.n1732 VSS.n1724 394
R1393 VSS.n1736 VSS.n1734 394
R1394 VSS.n1740 VSS.n1722 394
R1395 VSS.n1744 VSS.n1742 394
R1396 VSS.n1748 VSS.n1720 394
R1397 VSS.n1752 VSS.n1750 394
R1398 VSS.n1756 VSS.n1718 394
R1399 VSS.n1760 VSS.n1758 394
R1400 VSS.n1764 VSS.n1716 394
R1401 VSS.n1768 VSS.n1766 394
R1402 VSS.n1779 VSS.n808 394
R1403 VSS.n892 VSS.n808 394
R1404 VSS.n892 VSS.n816 394
R1405 VSS.n1773 VSS.n816 394
R1406 VSS.n1773 VSS.n1772 394
R1407 VSS.n1772 VSS.n834 394
R1408 VSS.n2010 VSS.n834 394
R1409 VSS.n2010 VSS.n333 394
R1410 VSS.n2004 VSS.n333 394
R1411 VSS.n2004 VSS.n341 394
R1412 VSS.n2252 VSS.n341 394
R1413 VSS.n362 VSS.n361 394
R1414 VSS.n2291 VSS.n361 394
R1415 VSS.n2289 VSS.n2288 394
R1416 VSS.n2285 VSS.n2284 394
R1417 VSS.n2281 VSS.n2280 394
R1418 VSS.n2277 VSS.n2276 394
R1419 VSS.n2273 VSS.n2272 394
R1420 VSS.n2269 VSS.n2268 394
R1421 VSS.n2265 VSS.n2264 394
R1422 VSS.n2261 VSS.n2260 394
R1423 VSS.n2257 VSS.n2256 394
R1424 VSS.n1639 VSS.n957 394
R1425 VSS.n1639 VSS.n938 394
R1426 VSS.n1659 VSS.n938 394
R1427 VSS.n1659 VSS.n936 394
R1428 VSS.n1663 VSS.n936 394
R1429 VSS.n1663 VSS.n917 394
R1430 VSS.n1683 VSS.n917 394
R1431 VSS.n1683 VSS.n915 394
R1432 VSS.n1687 VSS.n915 394
R1433 VSS.n1687 VSS.n736 394
R1434 VSS.n2052 VSS.n736 394
R1435 VSS.n1635 VSS.n959 394
R1436 VSS.n1632 VSS.n1579 394
R1437 VSS.n1628 VSS.n1627 394
R1438 VSS.n1624 VSS.n1623 394
R1439 VSS.n1620 VSS.n1619 394
R1440 VSS.n1616 VSS.n1615 394
R1441 VSS.n1612 VSS.n1611 394
R1442 VSS.n1608 VSS.n1607 394
R1443 VSS.n1604 VSS.n1603 394
R1444 VSS.n1600 VSS.n1599 394
R1445 VSS.n1596 VSS.n1595 394
R1446 VSS.n1591 VSS.n955 394
R1447 VSS.n955 VSS.n947 394
R1448 VSS.n947 VSS.n940 394
R1449 VSS.n1585 VSS.n940 394
R1450 VSS.n1585 VSS.n934 394
R1451 VSS.n934 VSS.n926 394
R1452 VSS.n926 VSS.n919 394
R1453 VSS.n1580 VSS.n919 394
R1454 VSS.n1580 VSS.n914 394
R1455 VSS.n914 VSS.n732 394
R1456 VSS.n2054 VSS.n732 394
R1457 VSS.n2048 VSS.n740 394
R1458 VSS.n752 VSS.n740 394
R1459 VSS.n756 VSS.n755 394
R1460 VSS.n760 VSS.n759 394
R1461 VSS.n764 VSS.n763 394
R1462 VSS.n768 VSS.n767 394
R1463 VSS.n772 VSS.n771 394
R1464 VSS.n776 VSS.n775 394
R1465 VSS.n780 VSS.n779 394
R1466 VSS.n784 VSS.n783 394
R1467 VSS.n788 VSS.n751 394
R1468 VSS.n1152 VSS.n1051 394
R1469 VSS.n1152 VSS.n1044 394
R1470 VSS.n1160 VSS.n1044 394
R1471 VSS.n1160 VSS.n1042 394
R1472 VSS.n1164 VSS.n1042 394
R1473 VSS.n1164 VSS.n1035 394
R1474 VSS.n1180 VSS.n1035 394
R1475 VSS.n1180 VSS.n1033 394
R1476 VSS.n1184 VSS.n1033 394
R1477 VSS.n1184 VSS.n1025 394
R1478 VSS.n1432 VSS.n1025 394
R1479 VSS.n1432 VSS.n1022 394
R1480 VSS.n1437 VSS.n1022 394
R1481 VSS.n1437 VSS.n1023 394
R1482 VSS.n1023 VSS.n1007 394
R1483 VSS.n1494 VSS.n1007 394
R1484 VSS.n1494 VSS.n1004 394
R1485 VSS.n1499 VSS.n1004 394
R1486 VSS.n1499 VSS.n1005 394
R1487 VSS.n1005 VSS.n989 394
R1488 VSS.n1518 VSS.n989 394
R1489 VSS.n1518 VSS.n986 394
R1490 VSS.n1523 VSS.n986 394
R1491 VSS.n1523 VSS.n987 394
R1492 VSS.n987 VSS.n965 394
R1493 VSS.n1563 VSS.n965 394
R1494 VSS.n1563 VSS.n963 394
R1495 VSS.n1567 VSS.n963 394
R1496 VSS.n1567 VSS.n951 394
R1497 VSS.n1643 VSS.n951 394
R1498 VSS.n1643 VSS.n949 394
R1499 VSS.n1647 VSS.n949 394
R1500 VSS.n1647 VSS.n930 394
R1501 VSS.n1667 VSS.n930 394
R1502 VSS.n1667 VSS.n928 394
R1503 VSS.n1671 VSS.n928 394
R1504 VSS.n1671 VSS.n909 394
R1505 VSS.n1691 VSS.n909 394
R1506 VSS.n1691 VSS.n906 394
R1507 VSS.n1696 VSS.n906 394
R1508 VSS.n1696 VSS.n907 394
R1509 VSS.n907 VSS.n792 394
R1510 VSS.n2044 VSS.n792 394
R1511 VSS.n2044 VSS.n793 394
R1512 VSS.n2040 VSS.n793 394
R1513 VSS.n2040 VSS.n796 394
R1514 VSS.n822 VSS.n796 394
R1515 VSS.n823 VSS.n822 394
R1516 VSS.n823 VSS.n819 394
R1517 VSS.n2023 VSS.n819 394
R1518 VSS.n2023 VSS.n820 394
R1519 VSS.n2019 VSS.n820 394
R1520 VSS.n2019 VSS.n831 394
R1521 VSS.n831 VSS.n830 394
R1522 VSS.n830 VSS.n827 394
R1523 VSS.n827 VSS.n344 394
R1524 VSS.n2304 VSS.n344 394
R1525 VSS.n2304 VSS.n345 394
R1526 VSS.n2300 VSS.n345 394
R1527 VSS.n2300 VSS.n348 394
R1528 VSS.n2150 VSS.n348 394
R1529 VSS.n1148 VSS.n1053 394
R1530 VSS.n1145 VSS.n1072 394
R1531 VSS.n1141 VSS.n1140 394
R1532 VSS.n1137 VSS.n1136 394
R1533 VSS.n1133 VSS.n1132 394
R1534 VSS.n1129 VSS.n1128 394
R1535 VSS.n1125 VSS.n1124 394
R1536 VSS.n1121 VSS.n1120 394
R1537 VSS.n1117 VSS.n1116 394
R1538 VSS.n1113 VSS.n1112 394
R1539 VSS.n1109 VSS.n1108 394
R1540 VSS.n1105 VSS.n1104 394
R1541 VSS.n1101 VSS.n1100 394
R1542 VSS.n1097 VSS.n1096 394
R1543 VSS.n1093 VSS.n1092 394
R1544 VSS.n1089 VSS.n1088 394
R1545 VSS.n1085 VSS.n1084 394
R1546 VSS.n1081 VSS.n1080 394
R1547 VSS.n1077 VSS.n1076 394
R1548 VSS.n1154 VSS.n1047 394
R1549 VSS.n1154 VSS.n1045 394
R1550 VSS.n1158 VSS.n1045 394
R1551 VSS.n1158 VSS.n1040 394
R1552 VSS.n1166 VSS.n1040 394
R1553 VSS.n1166 VSS.n1037 394
R1554 VSS.n1178 VSS.n1037 394
R1555 VSS.n1178 VSS.n1038 394
R1556 VSS.n1038 VSS.n1032 394
R1557 VSS.n1173 VSS.n1032 394
R1558 VSS.n1173 VSS.n1027 394
R1559 VSS.n1170 VSS.n1027 394
R1560 VSS.n1170 VSS.n1021 394
R1561 VSS.n1021 VSS.n1012 394
R1562 VSS.n1448 VSS.n1012 394
R1563 VSS.n1448 VSS.n1009 394
R1564 VSS.n1490 VSS.n1009 394
R1565 VSS.n1490 VSS.n1002 394
R1566 VSS.n1486 VSS.n1002 394
R1567 VSS.n1486 VSS.n1485 394
R1568 VSS.n1485 VSS.n991 394
R1569 VSS.n1481 VSS.n991 394
R1570 VSS.n1481 VSS.n984 394
R1571 VSS.n1478 VSS.n984 394
R1572 VSS.n1478 VSS.n1477 394
R1573 VSS.n1477 VSS.n967 394
R1574 VSS.n1472 VSS.n967 394
R1575 VSS.n1472 VSS.n961 394
R1576 VSS.n1469 VSS.n961 394
R1577 VSS.n1469 VSS.n953 394
R1578 VSS.n1466 VSS.n953 394
R1579 VSS.n1466 VSS.n948 394
R1580 VSS.n948 VSS.n941 394
R1581 VSS.n941 VSS.n932 394
R1582 VSS.n1461 VSS.n932 394
R1583 VSS.n1461 VSS.n927 394
R1584 VSS.n927 VSS.n920 394
R1585 VSS.n920 VSS.n911 394
R1586 VSS.n1456 VSS.n911 394
R1587 VSS.n1456 VSS.n905 394
R1588 VSS.n1453 VSS.n905 394
R1589 VSS.n1453 VSS.n1452 394
R1590 VSS.n1452 VSS.n790 394
R1591 VSS.n1789 VSS.n790 394
R1592 VSS.n1789 VSS.n798 394
R1593 VSS.n1793 VSS.n798 394
R1594 VSS.n1794 VSS.n1793 394
R1595 VSS.n1794 VSS.n893 394
R1596 VSS.n1798 VSS.n893 394
R1597 VSS.n1798 VSS.n817 394
R1598 VSS.n1993 VSS.n817 394
R1599 VSS.n1993 VSS.n833 394
R1600 VSS.n835 VSS.n833 394
R1601 VSS.n1997 VSS.n835 394
R1602 VSS.n1997 VSS.n839 394
R1603 VSS.n2001 VSS.n839 394
R1604 VSS.n2001 VSS.n342 394
R1605 VSS.n2157 VSS.n342 394
R1606 VSS.n2157 VSS.n349 394
R1607 VSS.n2153 VSS.n349 394
R1608 VSS.n2153 VSS.n2152 394
R1609 VSS.n2146 VSS.n370 394
R1610 VSS.n390 VSS.n370 394
R1611 VSS.n394 VSS.n393 394
R1612 VSS.n398 VSS.n397 394
R1613 VSS.n402 VSS.n401 394
R1614 VSS.n406 VSS.n405 394
R1615 VSS.n410 VSS.n409 394
R1616 VSS.n414 VSS.n413 394
R1617 VSS.n418 VSS.n417 394
R1618 VSS.n422 VSS.n421 394
R1619 VSS.n426 VSS.n425 394
R1620 VSS.n429 VSS.n428 394
R1621 VSS.n535 VSS.n534 394
R1622 VSS.n539 VSS.n538 394
R1623 VSS.n543 VSS.n542 394
R1624 VSS.n547 VSS.n546 394
R1625 VSS.n551 VSS.n550 394
R1626 VSS.n555 VSS.n554 394
R1627 VSS.n560 VSS.n388 394
R1628 VSS.n252 VSS.n236 394
R1629 VSS.n252 VSS.n230 394
R1630 VSS.n260 VSS.n230 394
R1631 VSS.n260 VSS.n228 394
R1632 VSS.n264 VSS.n228 394
R1633 VSS.n264 VSS.n222 394
R1634 VSS.n272 VSS.n222 394
R1635 VSS.n272 VSS.n220 394
R1636 VSS.n276 VSS.n220 394
R1637 VSS.n276 VSS.n214 394
R1638 VSS.n284 VSS.n214 394
R1639 VSS.n284 VSS.n212 394
R1640 VSS.n288 VSS.n212 394
R1641 VSS.n288 VSS.n203 394
R1642 VSS.n2386 VSS.n203 394
R1643 VSS.n2386 VSS.n204 394
R1644 VSS.n295 VSS.n204 394
R1645 VSS.n296 VSS.n295 394
R1646 VSS.n297 VSS.n296 394
R1647 VSS.n2184 VSS.n297 394
R1648 VSS.n2184 VSS.n302 394
R1649 VSS.n303 VSS.n302 394
R1650 VSS.n304 VSS.n303 394
R1651 VSS.n2240 VSS.n304 394
R1652 VSS.n2180 VSS.n2179 394
R1653 VSS.n2235 VSS.n2179 394
R1654 VSS.n2233 VSS.n2232 394
R1655 VSS.n2229 VSS.n2228 394
R1656 VSS.n2225 VSS.n2224 394
R1657 VSS.n2221 VSS.n2220 394
R1658 VSS.n2217 VSS.n2216 394
R1659 VSS.n2213 VSS.n2212 394
R1660 VSS.n2209 VSS.n2208 394
R1661 VSS.n2205 VSS.n2204 394
R1662 VSS.n2201 VSS.n2200 394
R1663 VSS.n2197 VSS.n2196 394
R1664 VSS.n2193 VSS.n2192 394
R1665 VSS.n2189 VSS.n2165 394
R1666 VSS.n2244 VSS.n2159 394
R1667 VSS.n2314 VSS.n331 394
R1668 VSS.n2161 VSS.n331 394
R1669 VSS.n2161 VSS.n2158 394
R1670 VSS.n2248 VSS.n2158 394
R1671 VSS.n254 VSS.n234 394
R1672 VSS.n254 VSS.n232 394
R1673 VSS.n258 VSS.n232 394
R1674 VSS.n258 VSS.n226 394
R1675 VSS.n266 VSS.n226 394
R1676 VSS.n266 VSS.n224 394
R1677 VSS.n270 VSS.n224 394
R1678 VSS.n270 VSS.n218 394
R1679 VSS.n278 VSS.n218 394
R1680 VSS.n278 VSS.n216 394
R1681 VSS.n282 VSS.n216 394
R1682 VSS.n282 VSS.n210 394
R1683 VSS.n290 VSS.n210 394
R1684 VSS.n290 VSS.n207 394
R1685 VSS.n2384 VSS.n207 394
R1686 VSS.n2384 VSS.n208 394
R1687 VSS.n2380 VSS.n208 394
R1688 VSS.n2380 VSS.n294 394
R1689 VSS.n2376 VSS.n294 394
R1690 VSS.n2376 VSS.n299 394
R1691 VSS.n2372 VSS.n299 394
R1692 VSS.n2372 VSS.n301 394
R1693 VSS.n2368 VSS.n301 394
R1694 VSS.n2368 VSS.n306 394
R1695 VSS.n2364 VSS.n2363 394
R1696 VSS.n2361 VSS.n310 394
R1697 VSS.n2357 VSS.n2356 394
R1698 VSS.n2354 VSS.n313 394
R1699 VSS.n2350 VSS.n2349 394
R1700 VSS.n2347 VSS.n316 394
R1701 VSS.n2343 VSS.n2342 394
R1702 VSS.n2340 VSS.n319 394
R1703 VSS.n2336 VSS.n2335 394
R1704 VSS.n2333 VSS.n322 394
R1705 VSS.n2329 VSS.n2328 394
R1706 VSS.n2326 VSS.n325 394
R1707 VSS.n2322 VSS.n2321 394
R1708 VSS.n2319 VSS.n328 394
R1709 VSS.n245 VSS.n240 394
R1710 VSS.n241 VSS.n238 394
R1711 VSS.n1440 VSS.n1018 394
R1712 VSS.n1440 VSS.n1015 394
R1713 VSS.n1445 VSS.n1015 394
R1714 VSS.n1445 VSS.n1016 394
R1715 VSS.n1016 VSS.n1000 394
R1716 VSS.n1502 VSS.n1000 394
R1717 VSS.n1502 VSS.n997 394
R1718 VSS.n1507 VSS.n997 394
R1719 VSS.n1507 VSS.n998 394
R1720 VSS.n998 VSS.n981 394
R1721 VSS.n1526 VSS.n981 394
R1722 VSS.n1526 VSS.n979 394
R1723 VSS.n1530 VSS.n979 394
R1724 VSS.n1530 VSS.n970 394
R1725 VSS.n1560 VSS.n970 394
R1726 VSS.n1560 VSS.n971 394
R1727 VSS.n1556 VSS.n971 394
R1728 VSS.n1556 VSS.n1555 394
R1729 VSS.n1555 VSS.n945 394
R1730 VSS.n1651 VSS.n945 394
R1731 VSS.n1651 VSS.n943 394
R1732 VSS.n1655 VSS.n943 394
R1733 VSS.n1655 VSS.n924 394
R1734 VSS.n1675 VSS.n924 394
R1735 VSS.n1675 VSS.n922 394
R1736 VSS.n1679 VSS.n922 394
R1737 VSS.n1679 VSS.n902 394
R1738 VSS.n1700 VSS.n902 394
R1739 VSS.n1700 VSS.n899 394
R1740 VSS.n1707 VSS.n899 394
R1741 VSS.n1707 VSS.n900 394
R1742 VSS.n1703 VSS.n900 394
R1743 VSS.n1703 VSS.n801 394
R1744 VSS.n2037 VSS.n801 394
R1745 VSS.n2037 VSS.n802 394
R1746 VSS.n2033 VSS.n802 394
R1747 VSS.n2033 VSS.n805 394
R1748 VSS.n889 VSS.n805 394
R1749 VSS.n888 VSS.n887 394
R1750 VSS.n1984 VSS.n887 394
R1751 VSS.n1982 VSS.n1981 394
R1752 VSS.n1978 VSS.n1977 394
R1753 VSS.n1974 VSS.n1973 394
R1754 VSS.n1970 VSS.n1969 394
R1755 VSS.n1966 VSS.n1965 394
R1756 VSS.n1962 VSS.n1961 394
R1757 VSS.n1958 VSS.n1957 394
R1758 VSS.n1954 VSS.n1953 394
R1759 VSS.n1950 VSS.n1949 394
R1760 VSS.n1942 VSS.n1941 394
R1761 VSS.n1938 VSS.n1937 394
R1762 VSS.n1934 VSS.n1933 394
R1763 VSS.n1930 VSS.n1929 394
R1764 VSS.n1926 VSS.n1925 394
R1765 VSS.n1922 VSS.n1921 394
R1766 VSS.n1918 VSS.n1917 394
R1767 VSS.n1914 VSS.n1913 394
R1768 VSS.n1910 VSS.n1909 394
R1769 VSS.n1906 VSS.n1905 394
R1770 VSS.n1902 VSS.n1901 394
R1771 VSS.n1894 VSS.n1893 394
R1772 VSS.n1890 VSS.n1889 394
R1773 VSS.n1886 VSS.n1885 394
R1774 VSS.n1882 VSS.n1881 394
R1775 VSS.n1878 VSS.n1877 394
R1776 VSS.n1874 VSS.n1873 394
R1777 VSS.n1870 VSS.n1869 394
R1778 VSS.n1866 VSS.n1865 394
R1779 VSS.n1862 VSS.n1861 394
R1780 VSS.n1858 VSS.n1857 394
R1781 VSS.n1854 VSS.n1853 394
R1782 VSS.n1846 VSS.n1845 394
R1783 VSS.n1842 VSS.n1841 394
R1784 VSS.n1838 VSS.n1837 394
R1785 VSS.n1834 VSS.n1833 394
R1786 VSS.n1830 VSS.n1829 394
R1787 VSS.n1826 VSS.n1825 394
R1788 VSS.n1822 VSS.n1821 394
R1789 VSS.n1818 VSS.n1817 394
R1790 VSS.n1814 VSS.n1813 394
R1791 VSS.n1810 VSS.n1809 394
R1792 VSS.n1806 VSS.n886 394
R1793 VSS.n1429 VSS.n1020 394
R1794 VSS.n1425 VSS.n1020 394
R1795 VSS.n1425 VSS.n1014 394
R1796 VSS.n1421 VSS.n1014 394
R1797 VSS.n1421 VSS.n1010 394
R1798 VSS.n1010 VSS.n1001 394
R1799 VSS.n1001 VSS.n994 394
R1800 VSS.n1509 VSS.n994 394
R1801 VSS.n1509 VSS.n992 394
R1802 VSS.n1515 VSS.n992 394
R1803 VSS.n1515 VSS.n983 394
R1804 VSS.n983 VSS.n977 394
R1805 VSS.n1532 VSS.n977 394
R1806 VSS.n1533 VSS.n1532 394
R1807 VSS.n1533 VSS.n968 394
R1808 VSS.n1536 VSS.n968 394
R1809 VSS.n1536 VSS.n975 394
R1810 VSS.n1553 VSS.n975 394
R1811 VSS.n1553 VSS.n954 394
R1812 VSS.n954 VSS.n946 394
R1813 VSS.n1548 VSS.n946 394
R1814 VSS.n1548 VSS.n942 394
R1815 VSS.n942 VSS.n933 394
R1816 VSS.n933 VSS.n925 394
R1817 VSS.n1543 VSS.n925 394
R1818 VSS.n1543 VSS.n921 394
R1819 VSS.n921 VSS.n912 394
R1820 VSS.n912 VSS.n904 394
R1821 VSS.n904 VSS.n897 394
R1822 VSS.n1709 VSS.n897 394
R1823 VSS.n1710 VSS.n1709 394
R1824 VSS.n1710 VSS.n895 394
R1825 VSS.n1786 VSS.n895 394
R1826 VSS.n1786 VSS.n799 394
R1827 VSS.n1782 VSS.n799 394
R1828 VSS.n1782 VSS.n807 394
R1829 VSS.n1802 VSS.n807 394
R1830 VSS.n1803 VSS.n1802 394
R1831 VSS.n1236 VSS.n1235 394
R1832 VSS.n1240 VSS.n1239 394
R1833 VSS.n1244 VSS.n1243 394
R1834 VSS.n1248 VSS.n1247 394
R1835 VSS.n1252 VSS.n1251 394
R1836 VSS.n1256 VSS.n1255 394
R1837 VSS.n1260 VSS.n1259 394
R1838 VSS.n1264 VSS.n1263 394
R1839 VSS.n1268 VSS.n1267 394
R1840 VSS.n1272 VSS.n1271 394
R1841 VSS.n1276 VSS.n1275 394
R1842 VSS.n1280 VSS.n1279 394
R1843 VSS.n1284 VSS.n1283 394
R1844 VSS.n1288 VSS.n1287 394
R1845 VSS.n1292 VSS.n1291 394
R1846 VSS.n1296 VSS.n1295 394
R1847 VSS.n1300 VSS.n1299 394
R1848 VSS.n1304 VSS.n1303 394
R1849 VSS.n1308 VSS.n1307 394
R1850 VSS.n1312 VSS.n1311 394
R1851 VSS.n1316 VSS.n1315 394
R1852 VSS.n1320 VSS.n1319 394
R1853 VSS.n1324 VSS.n1323 394
R1854 VSS.n1328 VSS.n1327 394
R1855 VSS.n1332 VSS.n1331 394
R1856 VSS.n1336 VSS.n1335 394
R1857 VSS.n1340 VSS.n1339 394
R1858 VSS.n1344 VSS.n1343 394
R1859 VSS.n1348 VSS.n1347 394
R1860 VSS.n1352 VSS.n1351 394
R1861 VSS.n1356 VSS.n1355 394
R1862 VSS.n1360 VSS.n1359 394
R1863 VSS.n1364 VSS.n1363 394
R1864 VSS.n1368 VSS.n1367 394
R1865 VSS.n1372 VSS.n1371 394
R1866 VSS.n1376 VSS.n1375 394
R1867 VSS.n1380 VSS.n1379 394
R1868 VSS.n1384 VSS.n1383 394
R1869 VSS.n1388 VSS.n1387 394
R1870 VSS.n1392 VSS.n1391 394
R1871 VSS.n1396 VSS.n1395 394
R1872 VSS.n1400 VSS.n1399 394
R1873 VSS.n1404 VSS.n1403 394
R1874 VSS.n1408 VSS.n1407 394
R1875 VSS.n1412 VSS.n1231 394
R1876 VSS.n1416 VSS.n1030 394
R1877 VSS.n724 VSS.n723 325.69
R1878 VSS.n669 VSS.n664 325.69
R1879 VSS.n1276 VSS.n1197 269.089
R1880 VSS.n1279 VSS.n1197 269.089
R1881 VSS.n191 VSS.t15 259.341
R1882 VSS.n108 VSS.t70 259.341
R1883 VSS.n91 VSS.t40 259.341
R1884 VSS.n8 VSS.t18 259.341
R1885 VSS.n190 VSS.t21 258.99
R1886 VSS.n189 VSS.t80 258.99
R1887 VSS.n188 VSS.t61 258.99
R1888 VSS.n101 VSS.t64 258.99
R1889 VSS.n102 VSS.t28 258.99
R1890 VSS.n105 VSS.t37 258.99
R1891 VSS.n106 VSS.t5 258.99
R1892 VSS.n107 VSS.t67 258.99
R1893 VSS.n90 VSS.t46 258.99
R1894 VSS.n89 VSS.t24 258.99
R1895 VSS.n88 VSS.t72 258.99
R1896 VSS.n1 VSS.t74 258.99
R1897 VSS.n2 VSS.t53 258.99
R1898 VSS.n5 VSS.t55 258.99
R1899 VSS.n6 VSS.t26 258.99
R1900 VSS.n7 VSS.t78 258.99
R1901 VSS.n183 VSS.n153 253.042
R1902 VSS.n123 VSS.n122 253.042
R1903 VSS.n86 VSS.n85 253.042
R1904 VSS.n22 VSS.n19 253.042
R1905 VSS.n246 VSS.n239 218.815
R1906 VSS.n247 VSS.n246 218.815
R1907 VSS.n2242 VSS.n2241 218.815
R1908 VSS.n2242 VSS.n2167 218.815
R1909 VSS.n2242 VSS.n2168 218.815
R1910 VSS.n2242 VSS.n2169 218.815
R1911 VSS.n2242 VSS.n2170 218.815
R1912 VSS.n2242 VSS.n2171 218.815
R1913 VSS.n2242 VSS.n2172 218.815
R1914 VSS.n2242 VSS.n2173 218.815
R1915 VSS.n2242 VSS.n2174 218.815
R1916 VSS.n2242 VSS.n2175 218.815
R1917 VSS.n2242 VSS.n2176 218.815
R1918 VSS.n2242 VSS.n2177 218.815
R1919 VSS.n2242 VSS.n2178 218.815
R1920 VSS.n2243 VSS.n2242 218.815
R1921 VSS.n330 VSS.n309 218.815
R1922 VSS.n2320 VSS.n309 218.815
R1923 VSS.n327 VSS.n309 218.815
R1924 VSS.n2327 VSS.n309 218.815
R1925 VSS.n324 VSS.n309 218.815
R1926 VSS.n2334 VSS.n309 218.815
R1927 VSS.n321 VSS.n309 218.815
R1928 VSS.n2341 VSS.n309 218.815
R1929 VSS.n318 VSS.n309 218.815
R1930 VSS.n2348 VSS.n309 218.815
R1931 VSS.n315 VSS.n309 218.815
R1932 VSS.n2355 VSS.n309 218.815
R1933 VSS.n312 VSS.n309 218.815
R1934 VSS.n2362 VSS.n309 218.815
R1935 VSS.n309 VSS.n308 218.815
R1936 VSS.n2145 VSS.n2144 218.815
R1937 VSS.n2144 VSS.n371 218.815
R1938 VSS.n2144 VSS.n372 218.815
R1939 VSS.n2144 VSS.n373 218.815
R1940 VSS.n2144 VSS.n374 218.815
R1941 VSS.n2144 VSS.n375 218.815
R1942 VSS.n2144 VSS.n376 218.815
R1943 VSS.n2144 VSS.n377 218.815
R1944 VSS.n2144 VSS.n378 218.815
R1945 VSS.n2144 VSS.n379 218.815
R1946 VSS.n2144 VSS.n380 218.815
R1947 VSS.n2144 VSS.n381 218.815
R1948 VSS.n2144 VSS.n382 218.815
R1949 VSS.n2144 VSS.n383 218.815
R1950 VSS.n2144 VSS.n384 218.815
R1951 VSS.n2144 VSS.n385 218.815
R1952 VSS.n2144 VSS.n386 218.815
R1953 VSS.n2144 VSS.n387 218.815
R1954 VSS.n2144 VSS.n561 218.815
R1955 VSS.n1147 VSS.n1054 218.815
R1956 VSS.n1147 VSS.n1055 218.815
R1957 VSS.n1147 VSS.n1056 218.815
R1958 VSS.n1147 VSS.n1057 218.815
R1959 VSS.n1147 VSS.n1058 218.815
R1960 VSS.n1147 VSS.n1059 218.815
R1961 VSS.n1147 VSS.n1060 218.815
R1962 VSS.n1147 VSS.n1061 218.815
R1963 VSS.n1147 VSS.n1062 218.815
R1964 VSS.n1147 VSS.n1063 218.815
R1965 VSS.n1147 VSS.n1064 218.815
R1966 VSS.n1147 VSS.n1065 218.815
R1967 VSS.n1147 VSS.n1066 218.815
R1968 VSS.n1147 VSS.n1067 218.815
R1969 VSS.n1147 VSS.n1068 218.815
R1970 VSS.n1147 VSS.n1069 218.815
R1971 VSS.n1147 VSS.n1070 218.815
R1972 VSS.n1147 VSS.n1071 218.815
R1973 VSS.n1147 VSS.n1146 218.815
R1974 VSS.n2047 VSS.n2046 218.815
R1975 VSS.n2046 VSS.n742 218.815
R1976 VSS.n2046 VSS.n743 218.815
R1977 VSS.n2046 VSS.n744 218.815
R1978 VSS.n2046 VSS.n745 218.815
R1979 VSS.n2046 VSS.n746 218.815
R1980 VSS.n2046 VSS.n747 218.815
R1981 VSS.n2046 VSS.n748 218.815
R1982 VSS.n2046 VSS.n749 218.815
R1983 VSS.n2046 VSS.n750 218.815
R1984 VSS.n2046 VSS.n789 218.815
R1985 VSS.n1634 VSS.n1569 218.815
R1986 VSS.n1634 VSS.n1570 218.815
R1987 VSS.n1634 VSS.n1571 218.815
R1988 VSS.n1634 VSS.n1572 218.815
R1989 VSS.n1634 VSS.n1573 218.815
R1990 VSS.n1634 VSS.n1574 218.815
R1991 VSS.n1634 VSS.n1575 218.815
R1992 VSS.n1634 VSS.n1576 218.815
R1993 VSS.n1634 VSS.n1577 218.815
R1994 VSS.n1634 VSS.n1578 218.815
R1995 VSS.n1634 VSS.n1633 218.815
R1996 VSS.n2298 VSS.n2297 218.815
R1997 VSS.n2298 VSS.n350 218.815
R1998 VSS.n2298 VSS.n351 218.815
R1999 VSS.n2298 VSS.n352 218.815
R2000 VSS.n2298 VSS.n353 218.815
R2001 VSS.n2298 VSS.n354 218.815
R2002 VSS.n2298 VSS.n355 218.815
R2003 VSS.n2298 VSS.n356 218.815
R2004 VSS.n2298 VSS.n357 218.815
R2005 VSS.n2298 VSS.n358 218.815
R2006 VSS.n2298 VSS.n359 218.815
R2007 VSS.n1767 VSS.n797 218.815
R2008 VSS.n1765 VSS.n797 218.815
R2009 VSS.n1759 VSS.n797 218.815
R2010 VSS.n1757 VSS.n797 218.815
R2011 VSS.n1751 VSS.n797 218.815
R2012 VSS.n1749 VSS.n797 218.815
R2013 VSS.n1743 VSS.n797 218.815
R2014 VSS.n1741 VSS.n797 218.815
R2015 VSS.n1735 VSS.n797 218.815
R2016 VSS.n1733 VSS.n797 218.815
R2017 VSS.n1727 VSS.n797 218.815
R2018 VSS.n2119 VSS.n2118 218.815
R2019 VSS.n2119 VSS.n585 218.815
R2020 VSS.n2119 VSS.n586 218.815
R2021 VSS.n2119 VSS.n587 218.815
R2022 VSS.n2119 VSS.n588 218.815
R2023 VSS.n2119 VSS.n589 218.815
R2024 VSS.n2119 VSS.n590 218.815
R2025 VSS.n2119 VSS.n591 218.815
R2026 VSS.n2119 VSS.n592 218.815
R2027 VSS.n2119 VSS.n593 218.815
R2028 VSS.n2119 VSS.n594 218.815
R2029 VSS.n651 VSS.n367 218.815
R2030 VSS.n600 VSS.n367 218.815
R2031 VSS.n644 VSS.n367 218.815
R2032 VSS.n638 VSS.n367 218.815
R2033 VSS.n636 VSS.n367 218.815
R2034 VSS.n630 VSS.n367 218.815
R2035 VSS.n628 VSS.n367 218.815
R2036 VSS.n622 VSS.n367 218.815
R2037 VSS.n620 VSS.n367 218.815
R2038 VSS.n614 VSS.n367 218.815
R2039 VSS.n612 VSS.n367 218.815
R2040 VSS.n1415 VSS.n1414 218.815
R2041 VSS.n1414 VSS.n1413 218.815
R2042 VSS.n1414 VSS.n1230 218.815
R2043 VSS.n1414 VSS.n1229 218.815
R2044 VSS.n1414 VSS.n1228 218.815
R2045 VSS.n1414 VSS.n1227 218.815
R2046 VSS.n1414 VSS.n1226 218.815
R2047 VSS.n1414 VSS.n1225 218.815
R2048 VSS.n1414 VSS.n1224 218.815
R2049 VSS.n1414 VSS.n1223 218.815
R2050 VSS.n1414 VSS.n1222 218.815
R2051 VSS.n1414 VSS.n1220 218.815
R2052 VSS.n1414 VSS.n1219 218.815
R2053 VSS.n1414 VSS.n1218 218.815
R2054 VSS.n1414 VSS.n1217 218.815
R2055 VSS.n1414 VSS.n1216 218.815
R2056 VSS.n1414 VSS.n1215 218.815
R2057 VSS.n1414 VSS.n1214 218.815
R2058 VSS.n1414 VSS.n1213 218.815
R2059 VSS.n1414 VSS.n1212 218.815
R2060 VSS.n1414 VSS.n1211 218.815
R2061 VSS.n1414 VSS.n1210 218.815
R2062 VSS.n1414 VSS.n1208 218.815
R2063 VSS.n1414 VSS.n1207 218.815
R2064 VSS.n1414 VSS.n1206 218.815
R2065 VSS.n1414 VSS.n1205 218.815
R2066 VSS.n1414 VSS.n1204 218.815
R2067 VSS.n1414 VSS.n1203 218.815
R2068 VSS.n1414 VSS.n1202 218.815
R2069 VSS.n1414 VSS.n1201 218.815
R2070 VSS.n1414 VSS.n1200 218.815
R2071 VSS.n1414 VSS.n1199 218.815
R2072 VSS.n1414 VSS.n1198 218.815
R2073 VSS.n1414 VSS.n1196 218.815
R2074 VSS.n1414 VSS.n1195 218.815
R2075 VSS.n1414 VSS.n1194 218.815
R2076 VSS.n1414 VSS.n1193 218.815
R2077 VSS.n1414 VSS.n1192 218.815
R2078 VSS.n1414 VSS.n1191 218.815
R2079 VSS.n1414 VSS.n1190 218.815
R2080 VSS.n1414 VSS.n1189 218.815
R2081 VSS.n1414 VSS.n1188 218.815
R2082 VSS.n1414 VSS.n1187 218.815
R2083 VSS.n1414 VSS.n1186 218.815
R2084 VSS.n1991 VSS.n1990 218.815
R2085 VSS.n1991 VSS.n841 218.815
R2086 VSS.n1991 VSS.n842 218.815
R2087 VSS.n1991 VSS.n843 218.815
R2088 VSS.n1991 VSS.n844 218.815
R2089 VSS.n1991 VSS.n845 218.815
R2090 VSS.n1991 VSS.n846 218.815
R2091 VSS.n1991 VSS.n847 218.815
R2092 VSS.n1991 VSS.n848 218.815
R2093 VSS.n1991 VSS.n849 218.815
R2094 VSS.n1991 VSS.n850 218.815
R2095 VSS.n1991 VSS.n851 218.815
R2096 VSS.n1991 VSS.n852 218.815
R2097 VSS.n1991 VSS.n853 218.815
R2098 VSS.n1991 VSS.n854 218.815
R2099 VSS.n1991 VSS.n855 218.815
R2100 VSS.n1991 VSS.n856 218.815
R2101 VSS.n1991 VSS.n857 218.815
R2102 VSS.n1991 VSS.n858 218.815
R2103 VSS.n1991 VSS.n859 218.815
R2104 VSS.n1991 VSS.n860 218.815
R2105 VSS.n1991 VSS.n861 218.815
R2106 VSS.n1991 VSS.n862 218.815
R2107 VSS.n1991 VSS.n863 218.815
R2108 VSS.n1991 VSS.n864 218.815
R2109 VSS.n1991 VSS.n865 218.815
R2110 VSS.n1991 VSS.n866 218.815
R2111 VSS.n1991 VSS.n867 218.815
R2112 VSS.n1991 VSS.n868 218.815
R2113 VSS.n1991 VSS.n869 218.815
R2114 VSS.n1991 VSS.n870 218.815
R2115 VSS.n1991 VSS.n871 218.815
R2116 VSS.n1991 VSS.n872 218.815
R2117 VSS.n1991 VSS.n873 218.815
R2118 VSS.n1991 VSS.n874 218.815
R2119 VSS.n1991 VSS.n875 218.815
R2120 VSS.n1991 VSS.n876 218.815
R2121 VSS.n1991 VSS.n877 218.815
R2122 VSS.n1991 VSS.n878 218.815
R2123 VSS.n1991 VSS.n879 218.815
R2124 VSS.n1991 VSS.n880 218.815
R2125 VSS.n1991 VSS.n881 218.815
R2126 VSS.n1991 VSS.n882 218.815
R2127 VSS.n1991 VSS.n883 218.815
R2128 VSS.n1991 VSS.n884 218.815
R2129 VSS.n1991 VSS.n885 218.815
R2130 VSS.n1324 VSS.n1209 198.87
R2131 VSS.n1372 VSS.n1221 198.87
R2132 VSS.n1375 VSS.n1221 198.87
R2133 VSS.n1327 VSS.n1209 198.87
R2134 VSS.n1414 VSS.n1221 193.066
R2135 VSS.n1414 VSS.n1209 193.066
R2136 VSS.n184 VSS.n183 185
R2137 VSS.n182 VSS.n181 185
R2138 VSS.n157 VSS.n156 185
R2139 VSS.n176 VSS.n175 185
R2140 VSS.n174 VSS.n173 185
R2141 VSS.n161 VSS.n160 185
R2142 VSS.n168 VSS.n167 185
R2143 VSS.n166 VSS.n165 185
R2144 VSS.n124 VSS.n123 185
R2145 VSS.n118 VSS.n117 185
R2146 VSS.n130 VSS.n129 185
R2147 VSS.n132 VSS.n131 185
R2148 VSS.n114 VSS.n113 185
R2149 VSS.n139 VSS.n138 185
R2150 VSS.n141 VSS.n140 185
R2151 VSS.n143 VSS.n110 185
R2152 VSS.n527 VSS.n526 185
R2153 VSS.n526 VSS.n525 185
R2154 VSS.n517 VSS.n516 185
R2155 VSS.n517 VSS.n512 185
R2156 VSS.n504 VSS.n496 185
R2157 VSS.n504 VSS.n495 185
R2158 VSS.n505 VSS.n504 185
R2159 VSS.n453 VSS.n452 185
R2160 VSS.n457 VSS.n452 185
R2161 VSS.n467 VSS.n466 185
R2162 VSS.n466 VSS.n465 185
R2163 VSS.n443 VSS.n435 185
R2164 VSS.n443 VSS.n434 185
R2165 VSS.n444 VSS.n443 185
R2166 VSS.n723 VSS.n722 185
R2167 VSS.n700 VSS.n699 185
R2168 VSS.n717 VSS.n716 185
R2169 VSS.n711 VSS.n710 185
R2170 VSS.n711 VSS.n703 185
R2171 VSS.n683 VSS.n682 185
R2172 VSS.n682 VSS.n681 185
R2173 VSS.n669 VSS.n668 185
R2174 VSS.n671 VSS.n670 185
R2175 VSS.n673 VSS.n661 185
R2176 VSS.n64 VSS.n63 185
R2177 VSS.n69 VSS.n68 185
R2178 VSS.n71 VSS.n70 185
R2179 VSS.n60 VSS.n59 185
R2180 VSS.n77 VSS.n76 185
R2181 VSS.n79 VSS.n78 185
R2182 VSS.n56 VSS.n55 185
R2183 VSS.n85 VSS.n84 185
R2184 VSS.n44 VSS.n43 185
R2185 VSS.n12 VSS.n11 185
R2186 VSS.n38 VSS.n37 185
R2187 VSS.n36 VSS.n35 185
R2188 VSS.n16 VSS.n15 185
R2189 VSS.n30 VSS.n29 185
R2190 VSS.n28 VSS.n27 185
R2191 VSS.n20 VSS.n19 185
R2192 VSS.n164 VSS.t17 178.418
R2193 VSS.t71 VSS.n144 178.418
R2194 VSS.n65 VSS.t42 178.418
R2195 VSS.t20 VSS.n10 178.418
R2196 VSS.t45 VSS.n715 175.332
R2197 VSS.t60 VSS.n674 175.332
R2198 VSS.n1414 VSS.n1197 157.957
R2199 VSS.n613 VSS.n612 147.374
R2200 VSS.n614 VSS.n608 147.374
R2201 VSS.n621 VSS.n620 147.374
R2202 VSS.n622 VSS.n606 147.374
R2203 VSS.n629 VSS.n628 147.374
R2204 VSS.n630 VSS.n604 147.374
R2205 VSS.n637 VSS.n636 147.374
R2206 VSS.n638 VSS.n602 147.374
R2207 VSS.n645 VSS.n644 147.374
R2208 VSS.n649 VSS.n600 147.374
R2209 VSS.n652 VSS.n651 147.374
R2210 VSS.n2118 VSS.n2117 147.374
R2211 VSS.n2112 VSS.n585 147.374
R2212 VSS.n2109 VSS.n586 147.374
R2213 VSS.n2105 VSS.n587 147.374
R2214 VSS.n2101 VSS.n588 147.374
R2215 VSS.n2097 VSS.n589 147.374
R2216 VSS.n2093 VSS.n590 147.374
R2217 VSS.n2089 VSS.n591 147.374
R2218 VSS.n2085 VSS.n592 147.374
R2219 VSS.n2081 VSS.n593 147.374
R2220 VSS.n2077 VSS.n594 147.374
R2221 VSS.n1727 VSS.n1724 147.374
R2222 VSS.n1734 VSS.n1733 147.374
R2223 VSS.n1735 VSS.n1722 147.374
R2224 VSS.n1742 VSS.n1741 147.374
R2225 VSS.n1743 VSS.n1720 147.374
R2226 VSS.n1750 VSS.n1749 147.374
R2227 VSS.n1751 VSS.n1718 147.374
R2228 VSS.n1758 VSS.n1757 147.374
R2229 VSS.n1759 VSS.n1716 147.374
R2230 VSS.n1766 VSS.n1765 147.374
R2231 VSS.n1767 VSS.n1714 147.374
R2232 VSS.n2297 VSS.n2296 147.374
R2233 VSS.n2291 VSS.n350 147.374
R2234 VSS.n2288 VSS.n351 147.374
R2235 VSS.n2284 VSS.n352 147.374
R2236 VSS.n2280 VSS.n353 147.374
R2237 VSS.n2276 VSS.n354 147.374
R2238 VSS.n2272 VSS.n355 147.374
R2239 VSS.n2268 VSS.n356 147.374
R2240 VSS.n2264 VSS.n357 147.374
R2241 VSS.n2260 VSS.n358 147.374
R2242 VSS.n2256 VSS.n359 147.374
R2243 VSS.n1633 VSS.n1632 147.374
R2244 VSS.n1628 VSS.n1578 147.374
R2245 VSS.n1624 VSS.n1577 147.374
R2246 VSS.n1620 VSS.n1576 147.374
R2247 VSS.n1616 VSS.n1575 147.374
R2248 VSS.n1612 VSS.n1574 147.374
R2249 VSS.n1608 VSS.n1573 147.374
R2250 VSS.n1604 VSS.n1572 147.374
R2251 VSS.n1600 VSS.n1571 147.374
R2252 VSS.n1596 VSS.n1570 147.374
R2253 VSS.n1592 VSS.n1569 147.374
R2254 VSS.n2047 VSS.n737 147.374
R2255 VSS.n752 VSS.n742 147.374
R2256 VSS.n756 VSS.n743 147.374
R2257 VSS.n760 VSS.n744 147.374
R2258 VSS.n764 VSS.n745 147.374
R2259 VSS.n768 VSS.n746 147.374
R2260 VSS.n772 VSS.n747 147.374
R2261 VSS.n776 VSS.n748 147.374
R2262 VSS.n780 VSS.n749 147.374
R2263 VSS.n784 VSS.n750 147.374
R2264 VSS.n789 VSS.n788 147.374
R2265 VSS.n1146 VSS.n1145 147.374
R2266 VSS.n1141 VSS.n1071 147.374
R2267 VSS.n1137 VSS.n1070 147.374
R2268 VSS.n1133 VSS.n1069 147.374
R2269 VSS.n1129 VSS.n1068 147.374
R2270 VSS.n1125 VSS.n1067 147.374
R2271 VSS.n1121 VSS.n1066 147.374
R2272 VSS.n1117 VSS.n1065 147.374
R2273 VSS.n1113 VSS.n1064 147.374
R2274 VSS.n1109 VSS.n1063 147.374
R2275 VSS.n1105 VSS.n1062 147.374
R2276 VSS.n1101 VSS.n1061 147.374
R2277 VSS.n1097 VSS.n1060 147.374
R2278 VSS.n1093 VSS.n1059 147.374
R2279 VSS.n1089 VSS.n1058 147.374
R2280 VSS.n1085 VSS.n1057 147.374
R2281 VSS.n1081 VSS.n1056 147.374
R2282 VSS.n1077 VSS.n1055 147.374
R2283 VSS.n1073 VSS.n1054 147.374
R2284 VSS.n2145 VSS.n368 147.374
R2285 VSS.n390 VSS.n371 147.374
R2286 VSS.n394 VSS.n372 147.374
R2287 VSS.n398 VSS.n373 147.374
R2288 VSS.n402 VSS.n374 147.374
R2289 VSS.n406 VSS.n375 147.374
R2290 VSS.n410 VSS.n376 147.374
R2291 VSS.n414 VSS.n377 147.374
R2292 VSS.n418 VSS.n378 147.374
R2293 VSS.n422 VSS.n379 147.374
R2294 VSS.n426 VSS.n380 147.374
R2295 VSS.n428 VSS.n381 147.374
R2296 VSS.n535 VSS.n382 147.374
R2297 VSS.n539 VSS.n383 147.374
R2298 VSS.n543 VSS.n384 147.374
R2299 VSS.n547 VSS.n385 147.374
R2300 VSS.n551 VSS.n386 147.374
R2301 VSS.n555 VSS.n387 147.374
R2302 VSS.n561 VSS.n560 147.374
R2303 VSS.n2241 VSS.n2240 147.374
R2304 VSS.n2235 VSS.n2167 147.374
R2305 VSS.n2232 VSS.n2168 147.374
R2306 VSS.n2228 VSS.n2169 147.374
R2307 VSS.n2224 VSS.n2170 147.374
R2308 VSS.n2220 VSS.n2171 147.374
R2309 VSS.n2216 VSS.n2172 147.374
R2310 VSS.n2212 VSS.n2173 147.374
R2311 VSS.n2208 VSS.n2174 147.374
R2312 VSS.n2204 VSS.n2175 147.374
R2313 VSS.n2200 VSS.n2176 147.374
R2314 VSS.n2196 VSS.n2177 147.374
R2315 VSS.n2192 VSS.n2178 147.374
R2316 VSS.n2243 VSS.n2165 147.374
R2317 VSS.n2364 VSS.n308 147.374
R2318 VSS.n2362 VSS.n2361 147.374
R2319 VSS.n2357 VSS.n312 147.374
R2320 VSS.n2355 VSS.n2354 147.374
R2321 VSS.n2350 VSS.n315 147.374
R2322 VSS.n2348 VSS.n2347 147.374
R2323 VSS.n2343 VSS.n318 147.374
R2324 VSS.n2341 VSS.n2340 147.374
R2325 VSS.n2336 VSS.n321 147.374
R2326 VSS.n2334 VSS.n2333 147.374
R2327 VSS.n2329 VSS.n324 147.374
R2328 VSS.n2327 VSS.n2326 147.374
R2329 VSS.n2322 VSS.n327 147.374
R2330 VSS.n2320 VSS.n2319 147.374
R2331 VSS.n2315 VSS.n330 147.374
R2332 VSS.n240 VSS.n239 147.374
R2333 VSS.n247 VSS.n238 147.374
R2334 VSS.n241 VSS.n239 147.374
R2335 VSS.n248 VSS.n247 147.374
R2336 VSS.n2241 VSS.n2180 147.374
R2337 VSS.n2233 VSS.n2167 147.374
R2338 VSS.n2229 VSS.n2168 147.374
R2339 VSS.n2225 VSS.n2169 147.374
R2340 VSS.n2221 VSS.n2170 147.374
R2341 VSS.n2217 VSS.n2171 147.374
R2342 VSS.n2213 VSS.n2172 147.374
R2343 VSS.n2209 VSS.n2173 147.374
R2344 VSS.n2205 VSS.n2174 147.374
R2345 VSS.n2201 VSS.n2175 147.374
R2346 VSS.n2197 VSS.n2176 147.374
R2347 VSS.n2193 VSS.n2177 147.374
R2348 VSS.n2189 VSS.n2178 147.374
R2349 VSS.n2244 VSS.n2243 147.374
R2350 VSS.n330 VSS.n328 147.374
R2351 VSS.n2321 VSS.n2320 147.374
R2352 VSS.n327 VSS.n325 147.374
R2353 VSS.n2328 VSS.n2327 147.374
R2354 VSS.n324 VSS.n322 147.374
R2355 VSS.n2335 VSS.n2334 147.374
R2356 VSS.n321 VSS.n319 147.374
R2357 VSS.n2342 VSS.n2341 147.374
R2358 VSS.n318 VSS.n316 147.374
R2359 VSS.n2349 VSS.n2348 147.374
R2360 VSS.n315 VSS.n313 147.374
R2361 VSS.n2356 VSS.n2355 147.374
R2362 VSS.n312 VSS.n310 147.374
R2363 VSS.n2363 VSS.n2362 147.374
R2364 VSS.n308 VSS.n306 147.374
R2365 VSS.n2146 VSS.n2145 147.374
R2366 VSS.n393 VSS.n371 147.374
R2367 VSS.n397 VSS.n372 147.374
R2368 VSS.n401 VSS.n373 147.374
R2369 VSS.n405 VSS.n374 147.374
R2370 VSS.n409 VSS.n375 147.374
R2371 VSS.n413 VSS.n376 147.374
R2372 VSS.n417 VSS.n377 147.374
R2373 VSS.n421 VSS.n378 147.374
R2374 VSS.n425 VSS.n379 147.374
R2375 VSS.n429 VSS.n380 147.374
R2376 VSS.n534 VSS.n381 147.374
R2377 VSS.n538 VSS.n382 147.374
R2378 VSS.n542 VSS.n383 147.374
R2379 VSS.n546 VSS.n384 147.374
R2380 VSS.n550 VSS.n385 147.374
R2381 VSS.n554 VSS.n386 147.374
R2382 VSS.n388 VSS.n387 147.374
R2383 VSS.n561 VSS.n366 147.374
R2384 VSS.n1076 VSS.n1054 147.374
R2385 VSS.n1080 VSS.n1055 147.374
R2386 VSS.n1084 VSS.n1056 147.374
R2387 VSS.n1088 VSS.n1057 147.374
R2388 VSS.n1092 VSS.n1058 147.374
R2389 VSS.n1096 VSS.n1059 147.374
R2390 VSS.n1100 VSS.n1060 147.374
R2391 VSS.n1104 VSS.n1061 147.374
R2392 VSS.n1108 VSS.n1062 147.374
R2393 VSS.n1112 VSS.n1063 147.374
R2394 VSS.n1116 VSS.n1064 147.374
R2395 VSS.n1120 VSS.n1065 147.374
R2396 VSS.n1124 VSS.n1066 147.374
R2397 VSS.n1128 VSS.n1067 147.374
R2398 VSS.n1132 VSS.n1068 147.374
R2399 VSS.n1136 VSS.n1069 147.374
R2400 VSS.n1140 VSS.n1070 147.374
R2401 VSS.n1072 VSS.n1071 147.374
R2402 VSS.n1146 VSS.n1053 147.374
R2403 VSS.n2048 VSS.n2047 147.374
R2404 VSS.n755 VSS.n742 147.374
R2405 VSS.n759 VSS.n743 147.374
R2406 VSS.n763 VSS.n744 147.374
R2407 VSS.n767 VSS.n745 147.374
R2408 VSS.n771 VSS.n746 147.374
R2409 VSS.n775 VSS.n747 147.374
R2410 VSS.n779 VSS.n748 147.374
R2411 VSS.n783 VSS.n749 147.374
R2412 VSS.n751 VSS.n750 147.374
R2413 VSS.n789 VSS.n733 147.374
R2414 VSS.n1595 VSS.n1569 147.374
R2415 VSS.n1599 VSS.n1570 147.374
R2416 VSS.n1603 VSS.n1571 147.374
R2417 VSS.n1607 VSS.n1572 147.374
R2418 VSS.n1611 VSS.n1573 147.374
R2419 VSS.n1615 VSS.n1574 147.374
R2420 VSS.n1619 VSS.n1575 147.374
R2421 VSS.n1623 VSS.n1576 147.374
R2422 VSS.n1627 VSS.n1577 147.374
R2423 VSS.n1579 VSS.n1578 147.374
R2424 VSS.n1633 VSS.n959 147.374
R2425 VSS.n2297 VSS.n362 147.374
R2426 VSS.n2289 VSS.n350 147.374
R2427 VSS.n2285 VSS.n351 147.374
R2428 VSS.n2281 VSS.n352 147.374
R2429 VSS.n2277 VSS.n353 147.374
R2430 VSS.n2273 VSS.n354 147.374
R2431 VSS.n2269 VSS.n355 147.374
R2432 VSS.n2265 VSS.n356 147.374
R2433 VSS.n2261 VSS.n357 147.374
R2434 VSS.n2257 VSS.n358 147.374
R2435 VSS.n2253 VSS.n359 147.374
R2436 VSS.n1768 VSS.n1767 147.374
R2437 VSS.n1765 VSS.n1764 147.374
R2438 VSS.n1760 VSS.n1759 147.374
R2439 VSS.n1757 VSS.n1756 147.374
R2440 VSS.n1752 VSS.n1751 147.374
R2441 VSS.n1749 VSS.n1748 147.374
R2442 VSS.n1744 VSS.n1743 147.374
R2443 VSS.n1741 VSS.n1740 147.374
R2444 VSS.n1736 VSS.n1735 147.374
R2445 VSS.n1733 VSS.n1732 147.374
R2446 VSS.n1728 VSS.n1727 147.374
R2447 VSS.n2118 VSS.n596 147.374
R2448 VSS.n2110 VSS.n585 147.374
R2449 VSS.n2106 VSS.n586 147.374
R2450 VSS.n2102 VSS.n587 147.374
R2451 VSS.n2098 VSS.n588 147.374
R2452 VSS.n2094 VSS.n589 147.374
R2453 VSS.n2090 VSS.n590 147.374
R2454 VSS.n2086 VSS.n591 147.374
R2455 VSS.n2082 VSS.n592 147.374
R2456 VSS.n2078 VSS.n593 147.374
R2457 VSS.n2074 VSS.n594 147.374
R2458 VSS.n651 VSS.n650 147.374
R2459 VSS.n646 VSS.n600 147.374
R2460 VSS.n644 VSS.n643 147.374
R2461 VSS.n639 VSS.n638 147.374
R2462 VSS.n636 VSS.n635 147.374
R2463 VSS.n631 VSS.n630 147.374
R2464 VSS.n628 VSS.n627 147.374
R2465 VSS.n623 VSS.n622 147.374
R2466 VSS.n620 VSS.n619 147.374
R2467 VSS.n615 VSS.n614 147.374
R2468 VSS.n612 VSS.n611 147.374
R2469 VSS.n1990 VSS.n1989 147.374
R2470 VSS.n1984 VSS.n841 147.374
R2471 VSS.n1981 VSS.n842 147.374
R2472 VSS.n1977 VSS.n843 147.374
R2473 VSS.n1973 VSS.n844 147.374
R2474 VSS.n1969 VSS.n845 147.374
R2475 VSS.n1965 VSS.n846 147.374
R2476 VSS.n1961 VSS.n847 147.374
R2477 VSS.n1957 VSS.n848 147.374
R2478 VSS.n1953 VSS.n849 147.374
R2479 VSS.n1949 VSS.n850 147.374
R2480 VSS.n1945 VSS.n851 147.374
R2481 VSS.n1941 VSS.n852 147.374
R2482 VSS.n1937 VSS.n853 147.374
R2483 VSS.n1933 VSS.n854 147.374
R2484 VSS.n1929 VSS.n855 147.374
R2485 VSS.n1925 VSS.n856 147.374
R2486 VSS.n1921 VSS.n857 147.374
R2487 VSS.n1917 VSS.n858 147.374
R2488 VSS.n1913 VSS.n859 147.374
R2489 VSS.n1909 VSS.n860 147.374
R2490 VSS.n1905 VSS.n861 147.374
R2491 VSS.n1901 VSS.n862 147.374
R2492 VSS.n1897 VSS.n863 147.374
R2493 VSS.n1893 VSS.n864 147.374
R2494 VSS.n1889 VSS.n865 147.374
R2495 VSS.n1885 VSS.n866 147.374
R2496 VSS.n1881 VSS.n867 147.374
R2497 VSS.n1877 VSS.n868 147.374
R2498 VSS.n1873 VSS.n869 147.374
R2499 VSS.n1869 VSS.n870 147.374
R2500 VSS.n1865 VSS.n871 147.374
R2501 VSS.n1861 VSS.n872 147.374
R2502 VSS.n1857 VSS.n873 147.374
R2503 VSS.n1853 VSS.n874 147.374
R2504 VSS.n1849 VSS.n875 147.374
R2505 VSS.n1845 VSS.n876 147.374
R2506 VSS.n1841 VSS.n877 147.374
R2507 VSS.n1837 VSS.n878 147.374
R2508 VSS.n1833 VSS.n879 147.374
R2509 VSS.n1829 VSS.n880 147.374
R2510 VSS.n1825 VSS.n881 147.374
R2511 VSS.n1821 VSS.n882 147.374
R2512 VSS.n1817 VSS.n883 147.374
R2513 VSS.n1813 VSS.n884 147.374
R2514 VSS.n1809 VSS.n885 147.374
R2515 VSS.n1232 VSS.n1186 147.374
R2516 VSS.n1236 VSS.n1187 147.374
R2517 VSS.n1240 VSS.n1188 147.374
R2518 VSS.n1244 VSS.n1189 147.374
R2519 VSS.n1248 VSS.n1190 147.374
R2520 VSS.n1252 VSS.n1191 147.374
R2521 VSS.n1256 VSS.n1192 147.374
R2522 VSS.n1260 VSS.n1193 147.374
R2523 VSS.n1264 VSS.n1194 147.374
R2524 VSS.n1268 VSS.n1195 147.374
R2525 VSS.n1272 VSS.n1196 147.374
R2526 VSS.n1280 VSS.n1198 147.374
R2527 VSS.n1284 VSS.n1199 147.374
R2528 VSS.n1288 VSS.n1200 147.374
R2529 VSS.n1292 VSS.n1201 147.374
R2530 VSS.n1296 VSS.n1202 147.374
R2531 VSS.n1300 VSS.n1203 147.374
R2532 VSS.n1304 VSS.n1204 147.374
R2533 VSS.n1308 VSS.n1205 147.374
R2534 VSS.n1312 VSS.n1206 147.374
R2535 VSS.n1316 VSS.n1207 147.374
R2536 VSS.n1320 VSS.n1208 147.374
R2537 VSS.n1328 VSS.n1210 147.374
R2538 VSS.n1332 VSS.n1211 147.374
R2539 VSS.n1336 VSS.n1212 147.374
R2540 VSS.n1340 VSS.n1213 147.374
R2541 VSS.n1344 VSS.n1214 147.374
R2542 VSS.n1348 VSS.n1215 147.374
R2543 VSS.n1352 VSS.n1216 147.374
R2544 VSS.n1356 VSS.n1217 147.374
R2545 VSS.n1360 VSS.n1218 147.374
R2546 VSS.n1364 VSS.n1219 147.374
R2547 VSS.n1368 VSS.n1220 147.374
R2548 VSS.n1376 VSS.n1222 147.374
R2549 VSS.n1380 VSS.n1223 147.374
R2550 VSS.n1384 VSS.n1224 147.374
R2551 VSS.n1388 VSS.n1225 147.374
R2552 VSS.n1392 VSS.n1226 147.374
R2553 VSS.n1396 VSS.n1227 147.374
R2554 VSS.n1400 VSS.n1228 147.374
R2555 VSS.n1404 VSS.n1229 147.374
R2556 VSS.n1408 VSS.n1230 147.374
R2557 VSS.n1413 VSS.n1412 147.374
R2558 VSS.n1416 VSS.n1415 147.374
R2559 VSS.n1415 VSS.n1028 147.374
R2560 VSS.n1413 VSS.n1030 147.374
R2561 VSS.n1231 VSS.n1230 147.374
R2562 VSS.n1407 VSS.n1229 147.374
R2563 VSS.n1403 VSS.n1228 147.374
R2564 VSS.n1399 VSS.n1227 147.374
R2565 VSS.n1395 VSS.n1226 147.374
R2566 VSS.n1391 VSS.n1225 147.374
R2567 VSS.n1387 VSS.n1224 147.374
R2568 VSS.n1383 VSS.n1223 147.374
R2569 VSS.n1379 VSS.n1222 147.374
R2570 VSS.n1371 VSS.n1220 147.374
R2571 VSS.n1367 VSS.n1219 147.374
R2572 VSS.n1363 VSS.n1218 147.374
R2573 VSS.n1359 VSS.n1217 147.374
R2574 VSS.n1355 VSS.n1216 147.374
R2575 VSS.n1351 VSS.n1215 147.374
R2576 VSS.n1347 VSS.n1214 147.374
R2577 VSS.n1343 VSS.n1213 147.374
R2578 VSS.n1339 VSS.n1212 147.374
R2579 VSS.n1335 VSS.n1211 147.374
R2580 VSS.n1331 VSS.n1210 147.374
R2581 VSS.n1323 VSS.n1208 147.374
R2582 VSS.n1319 VSS.n1207 147.374
R2583 VSS.n1315 VSS.n1206 147.374
R2584 VSS.n1311 VSS.n1205 147.374
R2585 VSS.n1307 VSS.n1204 147.374
R2586 VSS.n1303 VSS.n1203 147.374
R2587 VSS.n1299 VSS.n1202 147.374
R2588 VSS.n1295 VSS.n1201 147.374
R2589 VSS.n1291 VSS.n1200 147.374
R2590 VSS.n1287 VSS.n1199 147.374
R2591 VSS.n1283 VSS.n1198 147.374
R2592 VSS.n1275 VSS.n1196 147.374
R2593 VSS.n1271 VSS.n1195 147.374
R2594 VSS.n1267 VSS.n1194 147.374
R2595 VSS.n1263 VSS.n1193 147.374
R2596 VSS.n1259 VSS.n1192 147.374
R2597 VSS.n1255 VSS.n1191 147.374
R2598 VSS.n1251 VSS.n1190 147.374
R2599 VSS.n1247 VSS.n1189 147.374
R2600 VSS.n1243 VSS.n1188 147.374
R2601 VSS.n1239 VSS.n1187 147.374
R2602 VSS.n1235 VSS.n1186 147.374
R2603 VSS.n1990 VSS.n888 147.374
R2604 VSS.n1982 VSS.n841 147.374
R2605 VSS.n1978 VSS.n842 147.374
R2606 VSS.n1974 VSS.n843 147.374
R2607 VSS.n1970 VSS.n844 147.374
R2608 VSS.n1966 VSS.n845 147.374
R2609 VSS.n1962 VSS.n846 147.374
R2610 VSS.n1958 VSS.n847 147.374
R2611 VSS.n1954 VSS.n848 147.374
R2612 VSS.n1950 VSS.n849 147.374
R2613 VSS.n1946 VSS.n850 147.374
R2614 VSS.n1942 VSS.n851 147.374
R2615 VSS.n1938 VSS.n852 147.374
R2616 VSS.n1934 VSS.n853 147.374
R2617 VSS.n1930 VSS.n854 147.374
R2618 VSS.n1926 VSS.n855 147.374
R2619 VSS.n1922 VSS.n856 147.374
R2620 VSS.n1918 VSS.n857 147.374
R2621 VSS.n1914 VSS.n858 147.374
R2622 VSS.n1910 VSS.n859 147.374
R2623 VSS.n1906 VSS.n860 147.374
R2624 VSS.n1902 VSS.n861 147.374
R2625 VSS.n1898 VSS.n862 147.374
R2626 VSS.n1894 VSS.n863 147.374
R2627 VSS.n1890 VSS.n864 147.374
R2628 VSS.n1886 VSS.n865 147.374
R2629 VSS.n1882 VSS.n866 147.374
R2630 VSS.n1878 VSS.n867 147.374
R2631 VSS.n1874 VSS.n868 147.374
R2632 VSS.n1870 VSS.n869 147.374
R2633 VSS.n1866 VSS.n870 147.374
R2634 VSS.n1862 VSS.n871 147.374
R2635 VSS.n1858 VSS.n872 147.374
R2636 VSS.n1854 VSS.n873 147.374
R2637 VSS.n1850 VSS.n874 147.374
R2638 VSS.n1846 VSS.n875 147.374
R2639 VSS.n1842 VSS.n876 147.374
R2640 VSS.n1838 VSS.n877 147.374
R2641 VSS.n1834 VSS.n878 147.374
R2642 VSS.n1830 VSS.n879 147.374
R2643 VSS.n1826 VSS.n880 147.374
R2644 VSS.n1822 VSS.n881 147.374
R2645 VSS.n1818 VSS.n882 147.374
R2646 VSS.n1814 VSS.n883 147.374
R2647 VSS.n1810 VSS.n884 147.374
R2648 VSS.n1806 VSS.n885 147.374
R2649 VSS.n2119 VSS.n305 144.722
R2650 VSS.n183 VSS.n182 140.69
R2651 VSS.n182 VSS.n156 140.69
R2652 VSS.n175 VSS.n156 140.69
R2653 VSS.n175 VSS.n174 140.69
R2654 VSS.n174 VSS.n160 140.69
R2655 VSS.n167 VSS.n160 140.69
R2656 VSS.n167 VSS.n166 140.69
R2657 VSS.n123 VSS.n117 140.69
R2658 VSS.n130 VSS.n117 140.69
R2659 VSS.n131 VSS.n130 140.69
R2660 VSS.n131 VSS.n113 140.69
R2661 VSS.n139 VSS.n113 140.69
R2662 VSS.n140 VSS.n139 140.69
R2663 VSS.n140 VSS.n110 140.69
R2664 VSS.n723 VSS.n699 140.69
R2665 VSS.n716 VSS.n699 140.69
R2666 VSS.n670 VSS.n669 140.69
R2667 VSS.n670 VSS.n661 140.69
R2668 VSS.n69 VSS.n63 140.69
R2669 VSS.n70 VSS.n69 140.69
R2670 VSS.n70 VSS.n59 140.69
R2671 VSS.n77 VSS.n59 140.69
R2672 VSS.n78 VSS.n77 140.69
R2673 VSS.n78 VSS.n55 140.69
R2674 VSS.n85 VSS.n55 140.69
R2675 VSS.n44 VSS.n11 140.69
R2676 VSS.n37 VSS.n11 140.69
R2677 VSS.n37 VSS.n36 140.69
R2678 VSS.n36 VSS.n15 140.69
R2679 VSS.n29 VSS.n15 140.69
R2680 VSS.n29 VSS.n28 140.69
R2681 VSS.n28 VSS.n19 140.69
R2682 VSS.n2166 VSS.n305 91.4784
R2683 VSS.n521 VSS.t33 90.6265
R2684 VSS.n497 VSS.t14 90.6265
R2685 VSS.t52 VSS.n450 90.6265
R2686 VSS.n436 VSS.t36 90.6265
R2687 VSS.n244 VSS.n233 85.8358
R2688 VSS.n250 VSS.n249 85.8358
R2689 VSS.n2316 VSS.n329 85.8358
R2690 VSS.n2247 VSS.n2246 85.8358
R2691 VSS.n2141 VSS.n566 82.4476
R2692 VSS.n654 VSS.n653 82.4476
R2693 VSS.n2116 VSS.n581 82.4476
R2694 VSS.n2075 VSS.n2073 82.4476
R2695 VSS.n1725 VSS.n812 82.4476
R2696 VSS.n1778 VSS.n1770 82.4476
R2697 VSS.n2295 VSS.n338 82.4476
R2698 VSS.n2254 VSS.n363 82.4476
R2699 VSS.n1637 VSS.n1636 82.4476
R2700 VSS.n1593 VSS.n1590 82.4476
R2701 VSS.n2051 VSS.n2050 82.4476
R2702 VSS.n2055 VSS.n731 82.4476
R2703 VSS.n521 VSS.t31 81.8918
R2704 VSS.n520 VSS.t76 81.8918
R2705 VSS.n497 VSS.t11 81.8918
R2706 VSS.n461 VSS.t48 81.8918
R2707 VSS.n450 VSS.t51 81.8918
R2708 VSS.n436 VSS.t34 81.8918
R2709 VSS.n701 VSS.t8 81.8918
R2710 VSS.n714 VSS.t43 81.8918
R2711 VSS.n660 VSS.t59 81.8918
R2712 VSS.n677 VSS.t57 81.8918
R2713 VSS.n1150 VSS.n1149 76.8005
R2714 VSS.n2149 VSS.n2148 76.8005
R2715 VSS.n1074 VSS.n1046 76.8005
R2716 VSS.n558 VSS.n365 76.8005
R2717 VSS.n1233 VSS.n1017 76.8005
R2718 VSS.n1428 VSS.n1418 76.8005
R2719 VSS.n1988 VSS.n890 76.8005
R2720 VSS.n1805 VSS.n1804 76.8005
R2721 VSS.n166 VSS.t17 70.3453
R2722 VSS.t71 VSS.n110 70.3453
R2723 VSS.n716 VSS.t45 70.3453
R2724 VSS.t60 VSS.n661 70.3453
R2725 VSS.t42 VSS.n63 70.3453
R2726 VSS.t20 VSS.n44 70.3453
R2727 VSS.n1278 VSS.n1277 64.7534
R2728 VSS.n1947 VSS.n1944 64.7534
R2729 VSS.n246 VSS.n235 61.7668
R2730 VSS.n2120 VSS.n2119 41.8676
R2731 VSS.n1326 VSS.n1325 39.1534
R2732 VSS.n1374 VSS.n1373 39.1534
R2733 VSS.n1899 VSS.n1896 39.1534
R2734 VSS.n1851 VSS.n1848 39.1534
R2735 VSS.n1147 VSS.n1048 34.2854
R2736 VSS.n253 VSS.n235 33.0722
R2737 VSS.n253 VSS.n231 33.0722
R2738 VSS.n259 VSS.n231 33.0722
R2739 VSS.n259 VSS.n227 33.0722
R2740 VSS.n265 VSS.n227 33.0722
R2741 VSS.n265 VSS.n223 33.0722
R2742 VSS.n271 VSS.n223 33.0722
R2743 VSS.n271 VSS.n219 33.0722
R2744 VSS.n277 VSS.n219 33.0722
R2745 VSS.n277 VSS.n215 33.0722
R2746 VSS.n283 VSS.n215 33.0722
R2747 VSS.n283 VSS.n211 33.0722
R2748 VSS.n289 VSS.n211 33.0722
R2749 VSS.n289 VSS.n205 33.0722
R2750 VSS.n2385 VSS.n205 33.0722
R2751 VSS.n2385 VSS.n206 33.0722
R2752 VSS.n2379 VSS.n206 33.0722
R2753 VSS.n2379 VSS.n2378 33.0722
R2754 VSS.n2378 VSS.n2377 33.0722
R2755 VSS.n2377 VSS.n298 33.0722
R2756 VSS.n2371 VSS.n298 33.0722
R2757 VSS.n2371 VSS.n2370 33.0722
R2758 VSS.n2370 VSS.n2369 33.0722
R2759 VSS.n504 VSS.n503 32.8962
R2760 VSS.n443 VSS.n442 32.8962
R2761 VSS.n2144 VSS.n2143 29.3404
R2762 VSS.n717 VSS.n715 28.3989
R2763 VSS.n674 VSS.n673 28.3989
R2764 VSS.n489 VSS.n488 27.9576
R2765 VSS.n485 VSS.n484 27.9576
R2766 VSS.n481 VSS.n480 27.9576
R2767 VSS.n477 VSS.n476 27.9576
R2768 VSS.n473 VSS.n472 27.9576
R2769 VSS.n491 VSS.n490 27.7293
R2770 VSS.n487 VSS.n486 27.7293
R2771 VSS.n483 VSS.n482 27.7293
R2772 VSS.n479 VSS.n478 27.7293
R2773 VSS.n475 VSS.n474 27.7293
R2774 VSS.n471 VSS.n470 27.7293
R2775 VSS.n695 VSS.n694 27.7293
R2776 VSS.n693 VSS.n692 27.7293
R2777 VSS.n691 VSS.n690 27.7293
R2778 VSS.n689 VSS.n688 27.7293
R2779 VSS.n687 VSS.n686 27.7293
R2780 VSS.n526 VSS.n509 27.5286
R2781 VSS.n518 VSS.n517 27.5286
R2782 VSS.n459 VSS.n452 27.5286
R2783 VSS.n466 VSS.n449 27.5286
R2784 VSS.n711 VSS.n702 27.5286
R2785 VSS.n682 VSS.n659 27.5286
R2786 VSS.n187 VSS.n153 25.6009
R2787 VSS.n122 VSS.n121 25.6009
R2788 VSS.n87 VSS.n86 25.6009
R2789 VSS.n22 VSS.n21 25.6009
R2790 VSS.n610 VSS.n566 25.6005
R2791 VSS.n610 VSS.n609 25.6005
R2792 VSS.n616 VSS.n609 25.6005
R2793 VSS.n617 VSS.n616 25.6005
R2794 VSS.n618 VSS.n617 25.6005
R2795 VSS.n618 VSS.n607 25.6005
R2796 VSS.n624 VSS.n607 25.6005
R2797 VSS.n625 VSS.n624 25.6005
R2798 VSS.n626 VSS.n625 25.6005
R2799 VSS.n626 VSS.n605 25.6005
R2800 VSS.n632 VSS.n605 25.6005
R2801 VSS.n633 VSS.n632 25.6005
R2802 VSS.n634 VSS.n633 25.6005
R2803 VSS.n634 VSS.n603 25.6005
R2804 VSS.n640 VSS.n603 25.6005
R2805 VSS.n641 VSS.n640 25.6005
R2806 VSS.n642 VSS.n641 25.6005
R2807 VSS.n642 VSS.n601 25.6005
R2808 VSS.n647 VSS.n601 25.6005
R2809 VSS.n648 VSS.n647 25.6005
R2810 VSS.n648 VSS.n599 25.6005
R2811 VSS.n653 VSS.n599 25.6005
R2812 VSS.n2141 VSS.n2140 25.6005
R2813 VSS.n2140 VSS.n2139 25.6005
R2814 VSS.n2139 VSS.n567 25.6005
R2815 VSS.n2133 VSS.n567 25.6005
R2816 VSS.n2133 VSS.n2132 25.6005
R2817 VSS.n2132 VSS.n2131 25.6005
R2818 VSS.n2131 VSS.n574 25.6005
R2819 VSS.n2125 VSS.n574 25.6005
R2820 VSS.n2125 VSS.n2124 25.6005
R2821 VSS.n2124 VSS.n2123 25.6005
R2822 VSS.n2123 VSS.n581 25.6005
R2823 VSS.n2116 VSS.n2115 25.6005
R2824 VSS.n2115 VSS.n2114 25.6005
R2825 VSS.n2114 VSS.n2113 25.6005
R2826 VSS.n2113 VSS.n2111 25.6005
R2827 VSS.n2111 VSS.n2108 25.6005
R2828 VSS.n2108 VSS.n2107 25.6005
R2829 VSS.n2107 VSS.n2104 25.6005
R2830 VSS.n2104 VSS.n2103 25.6005
R2831 VSS.n2103 VSS.n2100 25.6005
R2832 VSS.n2100 VSS.n2099 25.6005
R2833 VSS.n2099 VSS.n2096 25.6005
R2834 VSS.n2096 VSS.n2095 25.6005
R2835 VSS.n2095 VSS.n2092 25.6005
R2836 VSS.n2092 VSS.n2091 25.6005
R2837 VSS.n2091 VSS.n2088 25.6005
R2838 VSS.n2088 VSS.n2087 25.6005
R2839 VSS.n2087 VSS.n2084 25.6005
R2840 VSS.n2084 VSS.n2083 25.6005
R2841 VSS.n2083 VSS.n2080 25.6005
R2842 VSS.n2080 VSS.n2079 25.6005
R2843 VSS.n2079 VSS.n2076 25.6005
R2844 VSS.n2076 VSS.n2075 25.6005
R2845 VSS.n2063 VSS.n2062 25.6005
R2846 VSS.n2064 VSS.n2063 25.6005
R2847 VSS.n2066 VSS.n2064 25.6005
R2848 VSS.n2067 VSS.n2066 25.6005
R2849 VSS.n2068 VSS.n2067 25.6005
R2850 VSS.n2069 VSS.n2068 25.6005
R2851 VSS.n2071 VSS.n2069 25.6005
R2852 VSS.n2072 VSS.n2071 25.6005
R2853 VSS.n2073 VSS.n2072 25.6005
R2854 VSS.n1729 VSS.n1725 25.6005
R2855 VSS.n1730 VSS.n1729 25.6005
R2856 VSS.n1731 VSS.n1730 25.6005
R2857 VSS.n1731 VSS.n1723 25.6005
R2858 VSS.n1737 VSS.n1723 25.6005
R2859 VSS.n1738 VSS.n1737 25.6005
R2860 VSS.n1739 VSS.n1738 25.6005
R2861 VSS.n1739 VSS.n1721 25.6005
R2862 VSS.n1745 VSS.n1721 25.6005
R2863 VSS.n1746 VSS.n1745 25.6005
R2864 VSS.n1747 VSS.n1746 25.6005
R2865 VSS.n1747 VSS.n1719 25.6005
R2866 VSS.n1753 VSS.n1719 25.6005
R2867 VSS.n1754 VSS.n1753 25.6005
R2868 VSS.n1755 VSS.n1754 25.6005
R2869 VSS.n1755 VSS.n1717 25.6005
R2870 VSS.n1761 VSS.n1717 25.6005
R2871 VSS.n1762 VSS.n1761 25.6005
R2872 VSS.n1763 VSS.n1762 25.6005
R2873 VSS.n1763 VSS.n1715 25.6005
R2874 VSS.n1769 VSS.n1715 25.6005
R2875 VSS.n1770 VSS.n1769 25.6005
R2876 VSS.n2029 VSS.n812 25.6005
R2877 VSS.n2029 VSS.n2028 25.6005
R2878 VSS.n2028 VSS.n2027 25.6005
R2879 VSS.n2027 VSS.n813 25.6005
R2880 VSS.n2014 VSS.n813 25.6005
R2881 VSS.n2015 VSS.n2014 25.6005
R2882 VSS.n2015 VSS.n337 25.6005
R2883 VSS.n2310 VSS.n337 25.6005
R2884 VSS.n2310 VSS.n2309 25.6005
R2885 VSS.n2309 VSS.n2308 25.6005
R2886 VSS.n2308 VSS.n338 25.6005
R2887 VSS.n2295 VSS.n2294 25.6005
R2888 VSS.n2294 VSS.n2293 25.6005
R2889 VSS.n2293 VSS.n2292 25.6005
R2890 VSS.n2292 VSS.n2290 25.6005
R2891 VSS.n2290 VSS.n2287 25.6005
R2892 VSS.n2287 VSS.n2286 25.6005
R2893 VSS.n2286 VSS.n2283 25.6005
R2894 VSS.n2283 VSS.n2282 25.6005
R2895 VSS.n2282 VSS.n2279 25.6005
R2896 VSS.n2279 VSS.n2278 25.6005
R2897 VSS.n2278 VSS.n2275 25.6005
R2898 VSS.n2275 VSS.n2274 25.6005
R2899 VSS.n2274 VSS.n2271 25.6005
R2900 VSS.n2271 VSS.n2270 25.6005
R2901 VSS.n2270 VSS.n2267 25.6005
R2902 VSS.n2267 VSS.n2266 25.6005
R2903 VSS.n2266 VSS.n2263 25.6005
R2904 VSS.n2263 VSS.n2262 25.6005
R2905 VSS.n2262 VSS.n2259 25.6005
R2906 VSS.n2259 VSS.n2258 25.6005
R2907 VSS.n2258 VSS.n2255 25.6005
R2908 VSS.n2255 VSS.n2254 25.6005
R2909 VSS.n1778 VSS.n1777 25.6005
R2910 VSS.n1777 VSS.n1776 25.6005
R2911 VSS.n1776 VSS.n1775 25.6005
R2912 VSS.n1775 VSS.n1774 25.6005
R2913 VSS.n1774 VSS.n1771 25.6005
R2914 VSS.n1771 VSS.n836 25.6005
R2915 VSS.n2009 VSS.n836 25.6005
R2916 VSS.n2005 VSS.n837 25.6005
R2917 VSS.n837 VSS.n363 25.6005
R2918 VSS.n1636 VSS.n958 25.6005
R2919 VSS.n1631 VSS.n958 25.6005
R2920 VSS.n1631 VSS.n1630 25.6005
R2921 VSS.n1630 VSS.n1629 25.6005
R2922 VSS.n1629 VSS.n1626 25.6005
R2923 VSS.n1626 VSS.n1625 25.6005
R2924 VSS.n1625 VSS.n1622 25.6005
R2925 VSS.n1622 VSS.n1621 25.6005
R2926 VSS.n1621 VSS.n1618 25.6005
R2927 VSS.n1618 VSS.n1617 25.6005
R2928 VSS.n1617 VSS.n1614 25.6005
R2929 VSS.n1614 VSS.n1613 25.6005
R2930 VSS.n1613 VSS.n1610 25.6005
R2931 VSS.n1610 VSS.n1609 25.6005
R2932 VSS.n1609 VSS.n1606 25.6005
R2933 VSS.n1606 VSS.n1605 25.6005
R2934 VSS.n1605 VSS.n1602 25.6005
R2935 VSS.n1602 VSS.n1601 25.6005
R2936 VSS.n1601 VSS.n1598 25.6005
R2937 VSS.n1598 VSS.n1597 25.6005
R2938 VSS.n1597 VSS.n1594 25.6005
R2939 VSS.n1594 VSS.n1593 25.6005
R2940 VSS.n1638 VSS.n1637 25.6005
R2941 VSS.n1638 VSS.n937 25.6005
R2942 VSS.n1660 VSS.n937 25.6005
R2943 VSS.n1661 VSS.n1660 25.6005
R2944 VSS.n1662 VSS.n1661 25.6005
R2945 VSS.n1662 VSS.n916 25.6005
R2946 VSS.n1684 VSS.n916 25.6005
R2947 VSS.n1685 VSS.n1684 25.6005
R2948 VSS.n1686 VSS.n1685 25.6005
R2949 VSS.n1686 VSS.n738 25.6005
R2950 VSS.n2051 VSS.n738 25.6005
R2951 VSS.n2050 VSS.n2049 25.6005
R2952 VSS.n2049 VSS.n739 25.6005
R2953 VSS.n753 VSS.n739 25.6005
R2954 VSS.n754 VSS.n753 25.6005
R2955 VSS.n757 VSS.n754 25.6005
R2956 VSS.n758 VSS.n757 25.6005
R2957 VSS.n761 VSS.n758 25.6005
R2958 VSS.n762 VSS.n761 25.6005
R2959 VSS.n765 VSS.n762 25.6005
R2960 VSS.n766 VSS.n765 25.6005
R2961 VSS.n769 VSS.n766 25.6005
R2962 VSS.n770 VSS.n769 25.6005
R2963 VSS.n773 VSS.n770 25.6005
R2964 VSS.n774 VSS.n773 25.6005
R2965 VSS.n777 VSS.n774 25.6005
R2966 VSS.n778 VSS.n777 25.6005
R2967 VSS.n781 VSS.n778 25.6005
R2968 VSS.n782 VSS.n781 25.6005
R2969 VSS.n785 VSS.n782 25.6005
R2970 VSS.n786 VSS.n785 25.6005
R2971 VSS.n787 VSS.n786 25.6005
R2972 VSS.n787 VSS.n731 25.6005
R2973 VSS.n1590 VSS.n1589 25.6005
R2974 VSS.n1589 VSS.n1588 25.6005
R2975 VSS.n1588 VSS.n1587 25.6005
R2976 VSS.n1587 VSS.n1586 25.6005
R2977 VSS.n1586 VSS.n1584 25.6005
R2978 VSS.n1584 VSS.n1583 25.6005
R2979 VSS.n1583 VSS.n1582 25.6005
R2980 VSS.n1582 VSS.n1581 25.6005
R2981 VSS.n913 VSS.n730 25.6005
R2982 VSS.n1151 VSS.n1150 25.6005
R2983 VSS.n1151 VSS.n1043 25.6005
R2984 VSS.n1161 VSS.n1043 25.6005
R2985 VSS.n1162 VSS.n1161 25.6005
R2986 VSS.n1163 VSS.n1162 25.6005
R2987 VSS.n1163 VSS.n1034 25.6005
R2988 VSS.n1181 VSS.n1034 25.6005
R2989 VSS.n1182 VSS.n1181 25.6005
R2990 VSS.n1183 VSS.n1182 25.6005
R2991 VSS.n1183 VSS.n1024 25.6005
R2992 VSS.n1433 VSS.n1024 25.6005
R2993 VSS.n1434 VSS.n1433 25.6005
R2994 VSS.n1436 VSS.n1434 25.6005
R2995 VSS.n1436 VSS.n1435 25.6005
R2996 VSS.n1435 VSS.n1006 25.6005
R2997 VSS.n1495 VSS.n1006 25.6005
R2998 VSS.n1496 VSS.n1495 25.6005
R2999 VSS.n1498 VSS.n1496 25.6005
R3000 VSS.n1498 VSS.n1497 25.6005
R3001 VSS.n1497 VSS.n988 25.6005
R3002 VSS.n1519 VSS.n988 25.6005
R3003 VSS.n1520 VSS.n1519 25.6005
R3004 VSS.n1522 VSS.n1520 25.6005
R3005 VSS.n1522 VSS.n1521 25.6005
R3006 VSS.n1521 VSS.n964 25.6005
R3007 VSS.n1564 VSS.n964 25.6005
R3008 VSS.n1565 VSS.n1564 25.6005
R3009 VSS.n1566 VSS.n1565 25.6005
R3010 VSS.n1566 VSS.n950 25.6005
R3011 VSS.n1644 VSS.n950 25.6005
R3012 VSS.n1645 VSS.n1644 25.6005
R3013 VSS.n1646 VSS.n1645 25.6005
R3014 VSS.n1646 VSS.n929 25.6005
R3015 VSS.n1668 VSS.n929 25.6005
R3016 VSS.n1669 VSS.n1668 25.6005
R3017 VSS.n1670 VSS.n1669 25.6005
R3018 VSS.n1670 VSS.n908 25.6005
R3019 VSS.n1692 VSS.n908 25.6005
R3020 VSS.n1693 VSS.n1692 25.6005
R3021 VSS.n1695 VSS.n1693 25.6005
R3022 VSS.n1695 VSS.n1694 25.6005
R3023 VSS.n1694 VSS.n794 25.6005
R3024 VSS.n2043 VSS.n794 25.6005
R3025 VSS.n2043 VSS.n2042 25.6005
R3026 VSS.n2042 VSS.n2041 25.6005
R3027 VSS.n2041 VSS.n795 25.6005
R3028 VSS.n821 VSS.n795 25.6005
R3029 VSS.n824 VSS.n821 25.6005
R3030 VSS.n825 VSS.n824 25.6005
R3031 VSS.n2022 VSS.n825 25.6005
R3032 VSS.n2022 VSS.n2021 25.6005
R3033 VSS.n2021 VSS.n2020 25.6005
R3034 VSS.n2020 VSS.n826 25.6005
R3035 VSS.n829 VSS.n826 25.6005
R3036 VSS.n829 VSS.n828 25.6005
R3037 VSS.n828 VSS.n346 25.6005
R3038 VSS.n2303 VSS.n346 25.6005
R3039 VSS.n2303 VSS.n2302 25.6005
R3040 VSS.n2302 VSS.n2301 25.6005
R3041 VSS.n2301 VSS.n347 25.6005
R3042 VSS.n2149 VSS.n347 25.6005
R3043 VSS.n1149 VSS.n1052 25.6005
R3044 VSS.n1144 VSS.n1052 25.6005
R3045 VSS.n1144 VSS.n1143 25.6005
R3046 VSS.n1143 VSS.n1142 25.6005
R3047 VSS.n1142 VSS.n1139 25.6005
R3048 VSS.n1139 VSS.n1138 25.6005
R3049 VSS.n1138 VSS.n1135 25.6005
R3050 VSS.n1135 VSS.n1134 25.6005
R3051 VSS.n1134 VSS.n1131 25.6005
R3052 VSS.n1131 VSS.n1130 25.6005
R3053 VSS.n1130 VSS.n1127 25.6005
R3054 VSS.n1127 VSS.n1126 25.6005
R3055 VSS.n1126 VSS.n1123 25.6005
R3056 VSS.n1123 VSS.n1122 25.6005
R3057 VSS.n1122 VSS.n1119 25.6005
R3058 VSS.n1119 VSS.n1118 25.6005
R3059 VSS.n1118 VSS.n1115 25.6005
R3060 VSS.n1115 VSS.n1114 25.6005
R3061 VSS.n1114 VSS.n1111 25.6005
R3062 VSS.n1111 VSS.n1110 25.6005
R3063 VSS.n1110 VSS.n1107 25.6005
R3064 VSS.n1107 VSS.n1106 25.6005
R3065 VSS.n1106 VSS.n1103 25.6005
R3066 VSS.n1103 VSS.n1102 25.6005
R3067 VSS.n1102 VSS.n1099 25.6005
R3068 VSS.n1099 VSS.n1098 25.6005
R3069 VSS.n1098 VSS.n1095 25.6005
R3070 VSS.n1095 VSS.n1094 25.6005
R3071 VSS.n1094 VSS.n1091 25.6005
R3072 VSS.n1091 VSS.n1090 25.6005
R3073 VSS.n1090 VSS.n1087 25.6005
R3074 VSS.n1087 VSS.n1086 25.6005
R3075 VSS.n1086 VSS.n1083 25.6005
R3076 VSS.n1083 VSS.n1082 25.6005
R3077 VSS.n1082 VSS.n1079 25.6005
R3078 VSS.n1079 VSS.n1078 25.6005
R3079 VSS.n1078 VSS.n1075 25.6005
R3080 VSS.n1075 VSS.n1074 25.6005
R3081 VSS.n1155 VSS.n1046 25.6005
R3082 VSS.n1156 VSS.n1155 25.6005
R3083 VSS.n1157 VSS.n1156 25.6005
R3084 VSS.n1157 VSS.n1039 25.6005
R3085 VSS.n1167 VSS.n1039 25.6005
R3086 VSS.n1168 VSS.n1167 25.6005
R3087 VSS.n1177 VSS.n1168 25.6005
R3088 VSS.n1177 VSS.n1176 25.6005
R3089 VSS.n1176 VSS.n1175 25.6005
R3090 VSS.n1175 VSS.n1174 25.6005
R3091 VSS.n1174 VSS.n1172 25.6005
R3092 VSS.n1172 VSS.n1171 25.6005
R3093 VSS.n1171 VSS.n1169 25.6005
R3094 VSS.n1169 VSS.n1011 25.6005
R3095 VSS.n1449 VSS.n1011 25.6005
R3096 VSS.n1450 VSS.n1449 25.6005
R3097 VSS.n1489 VSS.n1450 25.6005
R3098 VSS.n1489 VSS.n1488 25.6005
R3099 VSS.n1488 VSS.n1487 25.6005
R3100 VSS.n1487 VSS.n1484 25.6005
R3101 VSS.n1484 VSS.n1483 25.6005
R3102 VSS.n1483 VSS.n1482 25.6005
R3103 VSS.n1482 VSS.n1480 25.6005
R3104 VSS.n1480 VSS.n1479 25.6005
R3105 VSS.n1479 VSS.n1475 25.6005
R3106 VSS.n1475 VSS.n1474 25.6005
R3107 VSS.n1474 VSS.n1473 25.6005
R3108 VSS.n1473 VSS.n1471 25.6005
R3109 VSS.n1471 VSS.n1470 25.6005
R3110 VSS.n1470 VSS.n1468 25.6005
R3111 VSS.n1468 VSS.n1467 25.6005
R3112 VSS.n1467 VSS.n1465 25.6005
R3113 VSS.n1465 VSS.n1464 25.6005
R3114 VSS.n1464 VSS.n1463 25.6005
R3115 VSS.n1463 VSS.n1462 25.6005
R3116 VSS.n1462 VSS.n1460 25.6005
R3117 VSS.n1460 VSS.n1459 25.6005
R3118 VSS.n1459 VSS.n1458 25.6005
R3119 VSS.n1458 VSS.n1457 25.6005
R3120 VSS.n1457 VSS.n1455 25.6005
R3121 VSS.n1455 VSS.n1454 25.6005
R3122 VSS.n1454 VSS.n1451 25.6005
R3123 VSS.n1451 VSS.n894 25.6005
R3124 VSS.n1790 VSS.n894 25.6005
R3125 VSS.n1791 VSS.n1790 25.6005
R3126 VSS.n1792 VSS.n1791 25.6005
R3127 VSS.n1795 VSS.n1792 25.6005
R3128 VSS.n1796 VSS.n1795 25.6005
R3129 VSS.n1797 VSS.n1796 25.6005
R3130 VSS.n1797 VSS.n840 25.6005
R3131 VSS.n1994 VSS.n840 25.6005
R3132 VSS.n1995 VSS.n1994 25.6005
R3133 VSS.n1996 VSS.n1995 25.6005
R3134 VSS.n1998 VSS.n1996 25.6005
R3135 VSS.n1999 VSS.n1998 25.6005
R3136 VSS.n2000 VSS.n1999 25.6005
R3137 VSS.n2000 VSS.n364 25.6005
R3138 VSS.n2156 VSS.n364 25.6005
R3139 VSS.n2156 VSS.n2155 25.6005
R3140 VSS.n2155 VSS.n2154 25.6005
R3141 VSS.n2154 VSS.n365 25.6005
R3142 VSS.n2148 VSS.n2147 25.6005
R3143 VSS.n2147 VSS.n369 25.6005
R3144 VSS.n391 VSS.n369 25.6005
R3145 VSS.n392 VSS.n391 25.6005
R3146 VSS.n395 VSS.n392 25.6005
R3147 VSS.n396 VSS.n395 25.6005
R3148 VSS.n399 VSS.n396 25.6005
R3149 VSS.n400 VSS.n399 25.6005
R3150 VSS.n403 VSS.n400 25.6005
R3151 VSS.n404 VSS.n403 25.6005
R3152 VSS.n407 VSS.n404 25.6005
R3153 VSS.n408 VSS.n407 25.6005
R3154 VSS.n411 VSS.n408 25.6005
R3155 VSS.n412 VSS.n411 25.6005
R3156 VSS.n415 VSS.n412 25.6005
R3157 VSS.n416 VSS.n415 25.6005
R3158 VSS.n419 VSS.n416 25.6005
R3159 VSS.n420 VSS.n419 25.6005
R3160 VSS.n423 VSS.n420 25.6005
R3161 VSS.n424 VSS.n423 25.6005
R3162 VSS.n427 VSS.n424 25.6005
R3163 VSS.n430 VSS.n427 25.6005
R3164 VSS.n533 VSS.n389 25.6005
R3165 VSS.n536 VSS.n533 25.6005
R3166 VSS.n537 VSS.n536 25.6005
R3167 VSS.n540 VSS.n537 25.6005
R3168 VSS.n541 VSS.n540 25.6005
R3169 VSS.n544 VSS.n541 25.6005
R3170 VSS.n545 VSS.n544 25.6005
R3171 VSS.n548 VSS.n545 25.6005
R3172 VSS.n549 VSS.n548 25.6005
R3173 VSS.n552 VSS.n549 25.6005
R3174 VSS.n553 VSS.n552 25.6005
R3175 VSS.n556 VSS.n553 25.6005
R3176 VSS.n557 VSS.n556 25.6005
R3177 VSS.n559 VSS.n557 25.6005
R3178 VSS.n559 VSS.n558 25.6005
R3179 VSS.n244 VSS.n243 25.6005
R3180 VSS.n243 VSS.n242 25.6005
R3181 VSS.n242 VSS.n237 25.6005
R3182 VSS.n249 VSS.n237 25.6005
R3183 VSS.n255 VSS.n233 25.6005
R3184 VSS.n256 VSS.n255 25.6005
R3185 VSS.n257 VSS.n256 25.6005
R3186 VSS.n257 VSS.n225 25.6005
R3187 VSS.n267 VSS.n225 25.6005
R3188 VSS.n268 VSS.n267 25.6005
R3189 VSS.n269 VSS.n268 25.6005
R3190 VSS.n269 VSS.n217 25.6005
R3191 VSS.n279 VSS.n217 25.6005
R3192 VSS.n280 VSS.n279 25.6005
R3193 VSS.n281 VSS.n280 25.6005
R3194 VSS.n281 VSS.n209 25.6005
R3195 VSS.n291 VSS.n209 25.6005
R3196 VSS.n292 VSS.n291 25.6005
R3197 VSS.n2383 VSS.n292 25.6005
R3198 VSS.n2383 VSS.n2382 25.6005
R3199 VSS.n2382 VSS.n2381 25.6005
R3200 VSS.n2381 VSS.n293 25.6005
R3201 VSS.n2375 VSS.n293 25.6005
R3202 VSS.n2375 VSS.n2374 25.6005
R3203 VSS.n2374 VSS.n2373 25.6005
R3204 VSS.n2373 VSS.n300 25.6005
R3205 VSS.n2367 VSS.n300 25.6005
R3206 VSS.n2367 VSS.n2366 25.6005
R3207 VSS.n2366 VSS.n2365 25.6005
R3208 VSS.n2365 VSS.n307 25.6005
R3209 VSS.n2360 VSS.n307 25.6005
R3210 VSS.n2360 VSS.n2359 25.6005
R3211 VSS.n2359 VSS.n2358 25.6005
R3212 VSS.n2358 VSS.n311 25.6005
R3213 VSS.n2353 VSS.n311 25.6005
R3214 VSS.n2353 VSS.n2352 25.6005
R3215 VSS.n2352 VSS.n2351 25.6005
R3216 VSS.n2351 VSS.n314 25.6005
R3217 VSS.n2346 VSS.n314 25.6005
R3218 VSS.n2346 VSS.n2345 25.6005
R3219 VSS.n2345 VSS.n2344 25.6005
R3220 VSS.n2344 VSS.n317 25.6005
R3221 VSS.n2339 VSS.n317 25.6005
R3222 VSS.n2339 VSS.n2338 25.6005
R3223 VSS.n2338 VSS.n2337 25.6005
R3224 VSS.n2337 VSS.n320 25.6005
R3225 VSS.n2332 VSS.n320 25.6005
R3226 VSS.n2332 VSS.n2331 25.6005
R3227 VSS.n2331 VSS.n2330 25.6005
R3228 VSS.n2330 VSS.n323 25.6005
R3229 VSS.n2325 VSS.n323 25.6005
R3230 VSS.n2325 VSS.n2324 25.6005
R3231 VSS.n2324 VSS.n2323 25.6005
R3232 VSS.n2323 VSS.n326 25.6005
R3233 VSS.n2318 VSS.n326 25.6005
R3234 VSS.n2318 VSS.n2317 25.6005
R3235 VSS.n2317 VSS.n2316 25.6005
R3236 VSS.n2160 VSS.n329 25.6005
R3237 VSS.n2162 VSS.n2160 25.6005
R3238 VSS.n2163 VSS.n2162 25.6005
R3239 VSS.n2247 VSS.n2163 25.6005
R3240 VSS.n251 VSS.n250 25.6005
R3241 VSS.n251 VSS.n229 25.6005
R3242 VSS.n261 VSS.n229 25.6005
R3243 VSS.n262 VSS.n261 25.6005
R3244 VSS.n263 VSS.n262 25.6005
R3245 VSS.n263 VSS.n221 25.6005
R3246 VSS.n273 VSS.n221 25.6005
R3247 VSS.n274 VSS.n273 25.6005
R3248 VSS.n275 VSS.n274 25.6005
R3249 VSS.n275 VSS.n213 25.6005
R3250 VSS.n285 VSS.n213 25.6005
R3251 VSS.n286 VSS.n285 25.6005
R3252 VSS.n287 VSS.n286 25.6005
R3253 VSS.n287 VSS.n201 25.6005
R3254 VSS.n2387 VSS.n202 25.6005
R3255 VSS.n2181 VSS.n202 25.6005
R3256 VSS.n2182 VSS.n2181 25.6005
R3257 VSS.n2183 VSS.n2182 25.6005
R3258 VSS.n2185 VSS.n2183 25.6005
R3259 VSS.n2186 VSS.n2185 25.6005
R3260 VSS.n2187 VSS.n2186 25.6005
R3261 VSS.n2188 VSS.n2187 25.6005
R3262 VSS.n2239 VSS.n2188 25.6005
R3263 VSS.n2239 VSS.n2238 25.6005
R3264 VSS.n2238 VSS.n2237 25.6005
R3265 VSS.n2237 VSS.n2236 25.6005
R3266 VSS.n2236 VSS.n2234 25.6005
R3267 VSS.n2234 VSS.n2231 25.6005
R3268 VSS.n2231 VSS.n2230 25.6005
R3269 VSS.n2230 VSS.n2227 25.6005
R3270 VSS.n2227 VSS.n2226 25.6005
R3271 VSS.n2226 VSS.n2223 25.6005
R3272 VSS.n2223 VSS.n2222 25.6005
R3273 VSS.n2222 VSS.n2219 25.6005
R3274 VSS.n2219 VSS.n2218 25.6005
R3275 VSS.n2218 VSS.n2215 25.6005
R3276 VSS.n2215 VSS.n2214 25.6005
R3277 VSS.n2214 VSS.n2211 25.6005
R3278 VSS.n2211 VSS.n2210 25.6005
R3279 VSS.n2210 VSS.n2207 25.6005
R3280 VSS.n2207 VSS.n2206 25.6005
R3281 VSS.n2206 VSS.n2203 25.6005
R3282 VSS.n2203 VSS.n2202 25.6005
R3283 VSS.n2202 VSS.n2199 25.6005
R3284 VSS.n2199 VSS.n2198 25.6005
R3285 VSS.n2198 VSS.n2195 25.6005
R3286 VSS.n2195 VSS.n2194 25.6005
R3287 VSS.n2194 VSS.n2191 25.6005
R3288 VSS.n2191 VSS.n2190 25.6005
R3289 VSS.n2190 VSS.n2164 25.6005
R3290 VSS.n2245 VSS.n2164 25.6005
R3291 VSS.n2246 VSS.n2245 25.6005
R3292 VSS.n1234 VSS.n1233 25.6005
R3293 VSS.n1237 VSS.n1234 25.6005
R3294 VSS.n1238 VSS.n1237 25.6005
R3295 VSS.n1241 VSS.n1238 25.6005
R3296 VSS.n1242 VSS.n1241 25.6005
R3297 VSS.n1245 VSS.n1242 25.6005
R3298 VSS.n1246 VSS.n1245 25.6005
R3299 VSS.n1249 VSS.n1246 25.6005
R3300 VSS.n1250 VSS.n1249 25.6005
R3301 VSS.n1253 VSS.n1250 25.6005
R3302 VSS.n1254 VSS.n1253 25.6005
R3303 VSS.n1257 VSS.n1254 25.6005
R3304 VSS.n1258 VSS.n1257 25.6005
R3305 VSS.n1261 VSS.n1258 25.6005
R3306 VSS.n1262 VSS.n1261 25.6005
R3307 VSS.n1265 VSS.n1262 25.6005
R3308 VSS.n1266 VSS.n1265 25.6005
R3309 VSS.n1269 VSS.n1266 25.6005
R3310 VSS.n1270 VSS.n1269 25.6005
R3311 VSS.n1273 VSS.n1270 25.6005
R3312 VSS.n1274 VSS.n1273 25.6005
R3313 VSS.n1277 VSS.n1274 25.6005
R3314 VSS.n1281 VSS.n1278 25.6005
R3315 VSS.n1282 VSS.n1281 25.6005
R3316 VSS.n1285 VSS.n1282 25.6005
R3317 VSS.n1286 VSS.n1285 25.6005
R3318 VSS.n1289 VSS.n1286 25.6005
R3319 VSS.n1290 VSS.n1289 25.6005
R3320 VSS.n1293 VSS.n1290 25.6005
R3321 VSS.n1294 VSS.n1293 25.6005
R3322 VSS.n1297 VSS.n1294 25.6005
R3323 VSS.n1298 VSS.n1297 25.6005
R3324 VSS.n1301 VSS.n1298 25.6005
R3325 VSS.n1302 VSS.n1301 25.6005
R3326 VSS.n1305 VSS.n1302 25.6005
R3327 VSS.n1306 VSS.n1305 25.6005
R3328 VSS.n1309 VSS.n1306 25.6005
R3329 VSS.n1310 VSS.n1309 25.6005
R3330 VSS.n1313 VSS.n1310 25.6005
R3331 VSS.n1314 VSS.n1313 25.6005
R3332 VSS.n1317 VSS.n1314 25.6005
R3333 VSS.n1318 VSS.n1317 25.6005
R3334 VSS.n1321 VSS.n1318 25.6005
R3335 VSS.n1322 VSS.n1321 25.6005
R3336 VSS.n1325 VSS.n1322 25.6005
R3337 VSS.n1329 VSS.n1326 25.6005
R3338 VSS.n1330 VSS.n1329 25.6005
R3339 VSS.n1333 VSS.n1330 25.6005
R3340 VSS.n1334 VSS.n1333 25.6005
R3341 VSS.n1337 VSS.n1334 25.6005
R3342 VSS.n1338 VSS.n1337 25.6005
R3343 VSS.n1341 VSS.n1338 25.6005
R3344 VSS.n1342 VSS.n1341 25.6005
R3345 VSS.n1345 VSS.n1342 25.6005
R3346 VSS.n1346 VSS.n1345 25.6005
R3347 VSS.n1349 VSS.n1346 25.6005
R3348 VSS.n1350 VSS.n1349 25.6005
R3349 VSS.n1353 VSS.n1350 25.6005
R3350 VSS.n1354 VSS.n1353 25.6005
R3351 VSS.n1357 VSS.n1354 25.6005
R3352 VSS.n1358 VSS.n1357 25.6005
R3353 VSS.n1361 VSS.n1358 25.6005
R3354 VSS.n1362 VSS.n1361 25.6005
R3355 VSS.n1365 VSS.n1362 25.6005
R3356 VSS.n1366 VSS.n1365 25.6005
R3357 VSS.n1369 VSS.n1366 25.6005
R3358 VSS.n1370 VSS.n1369 25.6005
R3359 VSS.n1373 VSS.n1370 25.6005
R3360 VSS.n1377 VSS.n1374 25.6005
R3361 VSS.n1378 VSS.n1377 25.6005
R3362 VSS.n1381 VSS.n1378 25.6005
R3363 VSS.n1382 VSS.n1381 25.6005
R3364 VSS.n1385 VSS.n1382 25.6005
R3365 VSS.n1386 VSS.n1385 25.6005
R3366 VSS.n1389 VSS.n1386 25.6005
R3367 VSS.n1390 VSS.n1389 25.6005
R3368 VSS.n1393 VSS.n1390 25.6005
R3369 VSS.n1394 VSS.n1393 25.6005
R3370 VSS.n1397 VSS.n1394 25.6005
R3371 VSS.n1398 VSS.n1397 25.6005
R3372 VSS.n1401 VSS.n1398 25.6005
R3373 VSS.n1402 VSS.n1401 25.6005
R3374 VSS.n1405 VSS.n1402 25.6005
R3375 VSS.n1406 VSS.n1405 25.6005
R3376 VSS.n1409 VSS.n1406 25.6005
R3377 VSS.n1410 VSS.n1409 25.6005
R3378 VSS.n1411 VSS.n1410 25.6005
R3379 VSS.n1411 VSS.n1029 25.6005
R3380 VSS.n1417 VSS.n1029 25.6005
R3381 VSS.n1418 VSS.n1417 25.6005
R3382 VSS.n1441 VSS.n1017 25.6005
R3383 VSS.n1442 VSS.n1441 25.6005
R3384 VSS.n1444 VSS.n1442 25.6005
R3385 VSS.n1444 VSS.n1443 25.6005
R3386 VSS.n1443 VSS.n999 25.6005
R3387 VSS.n1503 VSS.n999 25.6005
R3388 VSS.n1504 VSS.n1503 25.6005
R3389 VSS.n1506 VSS.n1504 25.6005
R3390 VSS.n1506 VSS.n1505 25.6005
R3391 VSS.n1505 VSS.n980 25.6005
R3392 VSS.n1527 VSS.n980 25.6005
R3393 VSS.n1528 VSS.n1527 25.6005
R3394 VSS.n1529 VSS.n1528 25.6005
R3395 VSS.n1529 VSS.n972 25.6005
R3396 VSS.n1559 VSS.n972 25.6005
R3397 VSS.n1559 VSS.n1558 25.6005
R3398 VSS.n1558 VSS.n1557 25.6005
R3399 VSS.n1557 VSS.n973 25.6005
R3400 VSS.n973 VSS.n944 25.6005
R3401 VSS.n1652 VSS.n944 25.6005
R3402 VSS.n1653 VSS.n1652 25.6005
R3403 VSS.n1654 VSS.n1653 25.6005
R3404 VSS.n1654 VSS.n923 25.6005
R3405 VSS.n1676 VSS.n923 25.6005
R3406 VSS.n1677 VSS.n1676 25.6005
R3407 VSS.n1678 VSS.n1677 25.6005
R3408 VSS.n1678 VSS.n901 25.6005
R3409 VSS.n1701 VSS.n901 25.6005
R3410 VSS.n1702 VSS.n1701 25.6005
R3411 VSS.n1706 VSS.n1702 25.6005
R3412 VSS.n1706 VSS.n1705 25.6005
R3413 VSS.n1705 VSS.n1704 25.6005
R3414 VSS.n1704 VSS.n803 25.6005
R3415 VSS.n2036 VSS.n803 25.6005
R3416 VSS.n2036 VSS.n2035 25.6005
R3417 VSS.n2035 VSS.n2034 25.6005
R3418 VSS.n2034 VSS.n804 25.6005
R3419 VSS.n890 VSS.n804 25.6005
R3420 VSS.n1988 VSS.n1987 25.6005
R3421 VSS.n1987 VSS.n1986 25.6005
R3422 VSS.n1986 VSS.n1985 25.6005
R3423 VSS.n1985 VSS.n1983 25.6005
R3424 VSS.n1983 VSS.n1980 25.6005
R3425 VSS.n1980 VSS.n1979 25.6005
R3426 VSS.n1979 VSS.n1976 25.6005
R3427 VSS.n1976 VSS.n1975 25.6005
R3428 VSS.n1975 VSS.n1972 25.6005
R3429 VSS.n1972 VSS.n1971 25.6005
R3430 VSS.n1971 VSS.n1968 25.6005
R3431 VSS.n1968 VSS.n1967 25.6005
R3432 VSS.n1967 VSS.n1964 25.6005
R3433 VSS.n1964 VSS.n1963 25.6005
R3434 VSS.n1963 VSS.n1960 25.6005
R3435 VSS.n1960 VSS.n1959 25.6005
R3436 VSS.n1959 VSS.n1956 25.6005
R3437 VSS.n1956 VSS.n1955 25.6005
R3438 VSS.n1955 VSS.n1952 25.6005
R3439 VSS.n1952 VSS.n1951 25.6005
R3440 VSS.n1951 VSS.n1948 25.6005
R3441 VSS.n1948 VSS.n1947 25.6005
R3442 VSS.n1944 VSS.n1943 25.6005
R3443 VSS.n1943 VSS.n1940 25.6005
R3444 VSS.n1940 VSS.n1939 25.6005
R3445 VSS.n1939 VSS.n1936 25.6005
R3446 VSS.n1936 VSS.n1935 25.6005
R3447 VSS.n1935 VSS.n1932 25.6005
R3448 VSS.n1932 VSS.n1931 25.6005
R3449 VSS.n1931 VSS.n1928 25.6005
R3450 VSS.n1928 VSS.n1927 25.6005
R3451 VSS.n1927 VSS.n1924 25.6005
R3452 VSS.n1924 VSS.n1923 25.6005
R3453 VSS.n1923 VSS.n1920 25.6005
R3454 VSS.n1920 VSS.n1919 25.6005
R3455 VSS.n1919 VSS.n1916 25.6005
R3456 VSS.n1916 VSS.n1915 25.6005
R3457 VSS.n1915 VSS.n1912 25.6005
R3458 VSS.n1912 VSS.n1911 25.6005
R3459 VSS.n1911 VSS.n1908 25.6005
R3460 VSS.n1908 VSS.n1907 25.6005
R3461 VSS.n1907 VSS.n1904 25.6005
R3462 VSS.n1904 VSS.n1903 25.6005
R3463 VSS.n1903 VSS.n1900 25.6005
R3464 VSS.n1900 VSS.n1899 25.6005
R3465 VSS.n1896 VSS.n1895 25.6005
R3466 VSS.n1895 VSS.n1892 25.6005
R3467 VSS.n1892 VSS.n1891 25.6005
R3468 VSS.n1891 VSS.n1888 25.6005
R3469 VSS.n1888 VSS.n1887 25.6005
R3470 VSS.n1887 VSS.n1884 25.6005
R3471 VSS.n1884 VSS.n1883 25.6005
R3472 VSS.n1883 VSS.n1880 25.6005
R3473 VSS.n1880 VSS.n1879 25.6005
R3474 VSS.n1879 VSS.n1876 25.6005
R3475 VSS.n1876 VSS.n1875 25.6005
R3476 VSS.n1875 VSS.n1872 25.6005
R3477 VSS.n1872 VSS.n1871 25.6005
R3478 VSS.n1871 VSS.n1868 25.6005
R3479 VSS.n1868 VSS.n1867 25.6005
R3480 VSS.n1867 VSS.n1864 25.6005
R3481 VSS.n1864 VSS.n1863 25.6005
R3482 VSS.n1863 VSS.n1860 25.6005
R3483 VSS.n1860 VSS.n1859 25.6005
R3484 VSS.n1859 VSS.n1856 25.6005
R3485 VSS.n1856 VSS.n1855 25.6005
R3486 VSS.n1855 VSS.n1852 25.6005
R3487 VSS.n1852 VSS.n1851 25.6005
R3488 VSS.n1848 VSS.n1847 25.6005
R3489 VSS.n1847 VSS.n1844 25.6005
R3490 VSS.n1844 VSS.n1843 25.6005
R3491 VSS.n1843 VSS.n1840 25.6005
R3492 VSS.n1840 VSS.n1839 25.6005
R3493 VSS.n1839 VSS.n1836 25.6005
R3494 VSS.n1836 VSS.n1835 25.6005
R3495 VSS.n1835 VSS.n1832 25.6005
R3496 VSS.n1832 VSS.n1831 25.6005
R3497 VSS.n1831 VSS.n1828 25.6005
R3498 VSS.n1828 VSS.n1827 25.6005
R3499 VSS.n1827 VSS.n1824 25.6005
R3500 VSS.n1824 VSS.n1823 25.6005
R3501 VSS.n1823 VSS.n1820 25.6005
R3502 VSS.n1820 VSS.n1819 25.6005
R3503 VSS.n1819 VSS.n1816 25.6005
R3504 VSS.n1816 VSS.n1815 25.6005
R3505 VSS.n1815 VSS.n1812 25.6005
R3506 VSS.n1812 VSS.n1811 25.6005
R3507 VSS.n1811 VSS.n1808 25.6005
R3508 VSS.n1808 VSS.n1807 25.6005
R3509 VSS.n1807 VSS.n1805 25.6005
R3510 VSS.n1428 VSS.n1427 25.6005
R3511 VSS.n1427 VSS.n1426 25.6005
R3512 VSS.n1426 VSS.n1423 25.6005
R3513 VSS.n1423 VSS.n1422 25.6005
R3514 VSS.n1422 VSS.n1420 25.6005
R3515 VSS.n1420 VSS.n1419 25.6005
R3516 VSS.n1419 VSS.n993 25.6005
R3517 VSS.n1510 VSS.n993 25.6005
R3518 VSS.n1511 VSS.n1510 25.6005
R3519 VSS.n1514 VSS.n1511 25.6005
R3520 VSS.n1514 VSS.n1513 25.6005
R3521 VSS.n1513 VSS.n1512 25.6005
R3522 VSS.n1512 VSS.n976 25.6005
R3523 VSS.n1534 VSS.n976 25.6005
R3524 VSS.n1535 VSS.n1534 25.6005
R3525 VSS.n1537 VSS.n1535 25.6005
R3526 VSS.n1538 VSS.n1537 25.6005
R3527 VSS.n1552 VSS.n1538 25.6005
R3528 VSS.n1552 VSS.n1551 25.6005
R3529 VSS.n1551 VSS.n1550 25.6005
R3530 VSS.n1550 VSS.n1549 25.6005
R3531 VSS.n1549 VSS.n1547 25.6005
R3532 VSS.n1547 VSS.n1546 25.6005
R3533 VSS.n1546 VSS.n1545 25.6005
R3534 VSS.n1545 VSS.n1544 25.6005
R3535 VSS.n1544 VSS.n1542 25.6005
R3536 VSS.n1542 VSS.n1541 25.6005
R3537 VSS.n1541 VSS.n1540 25.6005
R3538 VSS.n1540 VSS.n1539 25.6005
R3539 VSS.n1539 VSS.n896 25.6005
R3540 VSS.n1711 VSS.n896 25.6005
R3541 VSS.n1712 VSS.n1711 25.6005
R3542 VSS.n1785 VSS.n1712 25.6005
R3543 VSS.n1785 VSS.n1784 25.6005
R3544 VSS.n1784 VSS.n1783 25.6005
R3545 VSS.n1783 VSS.n1713 25.6005
R3546 VSS.n1713 VSS.n891 25.6005
R3547 VSS.n1804 VSS.n891 25.6005
R3548 VSS.n185 VSS.n184 24.8476
R3549 VSS.n124 VSS.n120 24.8476
R3550 VSS.n502 VSS.n496 24.8476
R3551 VSS.n441 VSS.n435 24.8476
R3552 VSS.n718 VSS.n700 24.8476
R3553 VSS.n672 VSS.n671 24.8476
R3554 VSS.n2056 VSS.n2055 24.8476
R3555 VSS.n84 VSS.n54 24.8476
R3556 VSS.n23 VSS.n20 24.8476
R3557 VSS.n713 VSS.n712 24.75
R3558 VSS.n676 VSS.n675 24.75
R3559 VSS.n524 VSS.n509 24.2609
R3560 VSS.n518 VSS.n511 24.2609
R3561 VSS.n459 VSS.n458 24.2609
R3562 VSS.n464 VSS.n449 24.2609
R3563 VSS.n706 VSS.n702 24.2609
R3564 VSS.n680 VSS.n659 24.2609
R3565 VSS.n181 VSS.n155 23.3417
R3566 VSS.n125 VSS.n118 23.3417
R3567 VSS.n525 VSS.n524 23.3417
R3568 VSS.n512 VSS.n511 23.3417
R3569 VSS.n499 VSS.n495 23.3417
R3570 VSS.n458 VSS.n457 23.3417
R3571 VSS.n465 VSS.n464 23.3417
R3572 VSS.n438 VSS.n434 23.3417
R3573 VSS.n722 VSS.n721 23.3417
R3574 VSS.n706 VSS.n703 23.3417
R3575 VSS.n681 VSS.n680 23.3417
R3576 VSS.n668 VSS.n663 23.3417
R3577 VSS.n83 VSS.n56 23.3417
R3578 VSS.n27 VSS.n26 23.3417
R3579 VSS.n503 VSS.n502 22.4252
R3580 VSS.n442 VSS.n441 22.4252
R3581 VSS.n1153 VSS.n1048 22.4175
R3582 VSS.n1153 VSS.n1050 22.4175
R3583 VSS.n1159 VSS.n1041 22.4175
R3584 VSS.n1165 VSS.n1041 22.4175
R3585 VSS.n1179 VSS.n1036 22.4175
R3586 VSS.n1179 VSS.n1031 22.4175
R3587 VSS.n1185 VSS.n1031 22.4175
R3588 VSS.n1431 VSS.n1026 22.4175
R3589 VSS.n2151 VSS.n360 22.4175
R3590 VSS.n2143 VSS.n563 22.4175
R3591 VSS.n2137 VSS.n2136 22.4175
R3592 VSS.n2136 VSS.n2135 22.4175
R3593 VSS.n2135 VSS.n572 22.4175
R3594 VSS.n2129 VSS.n2128 22.4175
R3595 VSS.n2128 VSS.n2127 22.4175
R3596 VSS.n2127 VSS.n579 22.4175
R3597 VSS.n2121 VSS.n2120 22.4175
R3598 VSS.n180 VSS.n157 21.8358
R3599 VSS.n129 VSS.n128 21.8358
R3600 VSS.n527 VSS.n508 21.8358
R3601 VSS.n516 VSS.n515 21.8358
R3602 VSS.n505 VSS.n494 21.8358
R3603 VSS.n456 VSS.n453 21.8358
R3604 VSS.n467 VSS.n448 21.8358
R3605 VSS.n444 VSS.n433 21.8358
R3606 VSS.n724 VSS.n698 21.8358
R3607 VSS.n710 VSS.n709 21.8358
R3608 VSS.n683 VSS.n658 21.8358
R3609 VSS.n667 VSS.n664 21.8358
R3610 VSS.n1581 VSS.n729 21.8358
R3611 VSS.n80 VSS.n79 21.8358
R3612 VSS.n30 VSS.n18 21.8358
R3613 VSS.n2151 VSS.n367 21.7582
R3614 VSS.n1159 VSS.t35 21.4285
R3615 VSS.n431 VSS.n430 21.0829
R3616 VSS.n177 VSS.n176 20.3299
R3617 VSS.n132 VSS.n116 20.3299
R3618 VSS.n76 VSS.n58 20.3299
R3619 VSS.n31 VSS.n16 20.3299
R3620 VSS.n173 VSS.n159 18.824
R3621 VSS.n133 VSS.n114 18.824
R3622 VSS.n75 VSS.n60 18.824
R3623 VSS.n35 VSS.n34 18.824
R3624 VSS.n1165 VSS.t49 18.7912
R3625 VSS.n2007 VSS.n2006 18.0711
R3626 VSS.n172 VSS.n161 17.3181
R3627 VSS.n138 VSS.n137 17.3181
R3628 VSS.n72 VSS.n71 17.3181
R3629 VSS.n38 VSS.n14 17.3181
R3630 VSS.n165 VSS.n164 17.1928
R3631 VSS.n144 VSS.n143 17.1928
R3632 VSS.n65 VSS.n64 17.1928
R3633 VSS.n43 VSS.n10 17.1928
R3634 VSS.n2061 VSS.n598 16.9417
R3635 VSS.n2024 VSS.n818 16.8133
R3636 VSS.n2012 VSS.n2011 16.8133
R3637 VSS.t128 VSS.n563 15.8243
R3638 VSS.n2121 VSS.t98 15.8243
R3639 VSS.n169 VSS.n168 15.8123
R3640 VSS.n141 VSS.n112 15.8123
R3641 VSS.n68 VSS.n62 15.8123
R3642 VSS.n39 VSS.n12 15.8123
R3643 VSS.n2389 VSS.n2388 15.553
R3644 VSS.n2166 VSS.t123 14.8954
R3645 VSS.n528 VSS.n527 14.5711
R3646 VSS.n516 VSS.n513 14.5711
R3647 VSS.n506 VSS.n505 14.5711
R3648 VSS.n454 VSS.n453 14.5711
R3649 VSS.n468 VSS.n467 14.5711
R3650 VSS.n445 VSS.n444 14.5711
R3651 VSS.n725 VSS.n724 14.5711
R3652 VSS.n710 VSS.n704 14.5711
R3653 VSS.n684 VSS.n683 14.5711
R3654 VSS.n664 VSS.n656 14.5711
R3655 VSS.n165 VSS.n163 14.3064
R3656 VSS.n143 VSS.n142 14.3064
R3657 VSS.n67 VSS.n64 14.3064
R3658 VSS.n43 VSS.n42 14.3064
R3659 VSS.t103 VSS.n1185 14.176
R3660 VSS.n2299 VSS.n2298 13.8463
R3661 VSS.n2009 VSS.n2008 13.5534
R3662 VSS.n655 VSS.n598 13.177
R3663 VSS.n2388 VSS.n201 12.8005
R3664 VSS.n2388 VSS.n2387 12.8005
R3665 VSS.n2144 VSS.n367 12.5277
R3666 VSS.n655 VSS.n654 12.424
R3667 VSS.n2008 VSS.n2007 12.0476
R3668 VSS.n168 VSS.n163 11.2946
R3669 VSS.n142 VSS.n141 11.2946
R3670 VSS.n68 VSS.n67 11.2946
R3671 VSS.n42 VSS.n12 11.2946
R3672 VSS.n1431 VSS.n1430 11.209
R3673 VSS.n1430 VSS.n1019 11.209
R3674 VSS.n1439 VSS.n1019 11.209
R3675 VSS.n1439 VSS.n1438 11.209
R3676 VSS.n1424 VSS.n1013 11.209
R3677 VSS.n1446 VSS.n1013 11.209
R3678 VSS.n1447 VSS.n1446 11.209
R3679 VSS.n1447 VSS.n1008 11.209
R3680 VSS.n1493 VSS.n1008 11.209
R3681 VSS.n1493 VSS.n1492 11.209
R3682 VSS.n1492 VSS.n1491 11.209
R3683 VSS.n1501 VSS.n1500 11.209
R3684 VSS.n1500 VSS.n1003 11.209
R3685 VSS.n1003 VSS.n995 11.209
R3686 VSS.n1508 VSS.n995 11.209
R3687 VSS.n1508 VSS.n996 11.209
R3688 VSS.n996 VSS.n990 11.209
R3689 VSS.n1517 VSS.n990 11.209
R3690 VSS.n1516 VSS.n982 11.209
R3691 VSS.n1525 VSS.n982 11.209
R3692 VSS.n1525 VSS.n1524 11.209
R3693 VSS.n1524 VSS.n985 11.209
R3694 VSS.n985 VSS.n978 11.209
R3695 VSS.n1531 VSS.n978 11.209
R3696 VSS.n1476 VSS.n966 11.209
R3697 VSS.n1562 VSS.n966 11.209
R3698 VSS.n1562 VSS.n1561 11.209
R3699 VSS.n1561 VSS.n969 11.209
R3700 VSS.n969 VSS.n960 11.209
R3701 VSS.n1568 VSS.n962 11.209
R3702 VSS.n1554 VSS.n974 11.209
R3703 VSS.n1642 VSS.n1641 11.209
R3704 VSS.n1657 VSS.n1656 11.209
R3705 VSS.n1666 VSS.n1665 11.209
R3706 VSS.n1681 VSS.n1680 11.209
R3707 VSS.n1690 VSS.n1689 11.209
R3708 VSS.n1699 VSS.n903 11.209
R3709 VSS.n1697 VSS.n734 11.209
R3710 VSS.n1708 VSS.n735 11.209
R3711 VSS.n1708 VSS.n898 11.209
R3712 VSS.n898 VSS.n741 11.209
R3713 VSS.n2045 VSS.n791 11.209
R3714 VSS.n1788 VSS.n1787 11.209
R3715 VSS.n2039 VSS.n2038 11.209
R3716 VSS.n2038 VSS.n800 11.209
R3717 VSS.n1781 VSS.n800 11.209
R3718 VSS.n2032 VSS.n806 11.209
R3719 VSS.n1799 VSS.n815 11.209
R3720 VSS.t126 VSS.n2017 11.209
R3721 VSS.t125 VSS.n572 11.209
R3722 VSS.n2129 VSS.t125 11.209
R3723 VSS.n93 VSS.n92 11.0636
R3724 VSS.n94 VSS.n52 11.0636
R3725 VSS.n95 VSS.n51 11.0636
R3726 VSS.n96 VSS.n4 11.0636
R3727 VSS.n45 VSS.n9 11.0636
R3728 VSS.n47 VSS.n46 11.0636
R3729 VSS.n49 VSS.n48 11.0636
R3730 VSS.n50 VSS.n3 11.0636
R3731 VSS.n98 VSS.n97 11.0636
R3732 VSS.n193 VSS.n192 11.0636
R3733 VSS.n194 VSS.n152 11.0636
R3734 VSS.n195 VSS.n151 11.0636
R3735 VSS.n196 VSS.n104 11.0636
R3736 VSS.n145 VSS.n109 11.0636
R3737 VSS.n147 VSS.n146 11.0636
R3738 VSS.n149 VSS.n148 11.0636
R3739 VSS.n150 VSS.n103 11.0636
R3740 VSS.n198 VSS.n197 11.0636
R3741 VSS.t6 VSS.n1516 10.8793
R3742 VSS.n2313 VSS.n332 10.8793
R3743 VSS.n2305 VSS.n343 10.8793
R3744 VSS.n2250 VSS.n2249 10.8793
R3745 VSS.n2046 VSS.n2045 10.5497
R3746 VSS.n2249 VSS.t12 10.5497
R3747 VSS.t124 VSS.n809 10.22
R3748 VSS.t3 VSS.n340 9.89036
R3749 VSS.n169 VSS.n161 9.78874
R3750 VSS.n138 VSS.n112 9.78874
R3751 VSS.n71 VSS.n62 9.78874
R3752 VSS.n39 VSS.n38 9.78874
R3753 VSS.n185 VSS.n153 9.58499
R3754 VSS.n122 VSS.n120 9.58499
R3755 VSS.n86 VSS.n54 9.58499
R3756 VSS.n23 VSS.n22 9.58499
R3757 VSS.n1438 VSS.t19 9.5607
R3758 VSS.n2060 VSS.n655 9.41955
R3759 VSS.n2008 VSS.n728 9.41955
R3760 VSS.n2057 VSS.n729 9.41955
R3761 VSS.n532 VSS.n431 9.40467
R3762 VSS.n186 VSS.n185 9.3005
R3763 VSS.n155 VSS.n154 9.3005
R3764 VSS.n180 VSS.n179 9.3005
R3765 VSS.n178 VSS.n177 9.3005
R3766 VSS.n159 VSS.n158 9.3005
R3767 VSS.n172 VSS.n171 9.3005
R3768 VSS.n170 VSS.n169 9.3005
R3769 VSS.n163 VSS.n162 9.3005
R3770 VSS.n120 VSS.n119 9.3005
R3771 VSS.n126 VSS.n125 9.3005
R3772 VSS.n128 VSS.n127 9.3005
R3773 VSS.n116 VSS.n115 9.3005
R3774 VSS.n134 VSS.n133 9.3005
R3775 VSS.n137 VSS.n136 9.3005
R3776 VSS.n135 VSS.n112 9.3005
R3777 VSS.n142 VSS.n111 9.3005
R3778 VSS.n511 VSS.n510 9.3005
R3779 VSS.n515 VSS.n514 9.3005
R3780 VSS.n502 VSS.n501 9.3005
R3781 VSS.n500 VSS.n499 9.3005
R3782 VSS.n494 VSS.n493 9.3005
R3783 VSS.n524 VSS.n523 9.3005
R3784 VSS.n508 VSS.n507 9.3005
R3785 VSS.n464 VSS.n463 9.3005
R3786 VSS.n448 VSS.n447 9.3005
R3787 VSS.n441 VSS.n440 9.3005
R3788 VSS.n439 VSS.n438 9.3005
R3789 VSS.n433 VSS.n432 9.3005
R3790 VSS.n458 VSS.n451 9.3005
R3791 VSS.n456 VSS.n455 9.3005
R3792 VSS.n707 VSS.n706 9.3005
R3793 VSS.n709 VSS.n708 9.3005
R3794 VSS.n719 VSS.n718 9.3005
R3795 VSS.n721 VSS.n720 9.3005
R3796 VSS.n698 VSS.n697 9.3005
R3797 VSS.n672 VSS.n662 9.3005
R3798 VSS.n665 VSS.n663 9.3005
R3799 VSS.n667 VSS.n666 9.3005
R3800 VSS.n680 VSS.n679 9.3005
R3801 VSS.n658 VSS.n657 9.3005
R3802 VSS.n2061 VSS.n2060 9.3005
R3803 VSS.n2006 VSS.n728 9.3005
R3804 VSS.n2057 VSS.n2056 9.3005
R3805 VSS.n533 VSS.n532 9.3005
R3806 VSS.n944 VSS.n200 9.3005
R3807 VSS.n54 VSS.n53 9.3005
R3808 VSS.n83 VSS.n82 9.3005
R3809 VSS.n81 VSS.n80 9.3005
R3810 VSS.n58 VSS.n57 9.3005
R3811 VSS.n75 VSS.n74 9.3005
R3812 VSS.n73 VSS.n72 9.3005
R3813 VSS.n62 VSS.n61 9.3005
R3814 VSS.n67 VSS.n66 9.3005
R3815 VSS.n24 VSS.n23 9.3005
R3816 VSS.n26 VSS.n25 9.3005
R3817 VSS.n18 VSS.n17 9.3005
R3818 VSS.n32 VSS.n31 9.3005
R3819 VSS.n34 VSS.n33 9.3005
R3820 VSS.n14 VSS.n13 9.3005
R3821 VSS.n40 VSS.n39 9.3005
R3822 VSS.n42 VSS.n41 9.3005
R3823 VSS.n1551 VSS.n100 9.3005
R3824 VSS.n974 VSS.t29 8.90138
R3825 VSS.n1648 VSS.t65 8.90138
R3826 VSS.n2062 VSS.n2061 8.65932
R3827 VSS.n1787 VSS.n797 8.57171
R3828 VSS.t106 VSS.n832 8.57171
R3829 VSS.n2298 VSS.n360 8.57171
R3830 VSS.n173 VSS.n172 8.28285
R3831 VSS.n137 VSS.n114 8.28285
R3832 VSS.n72 VSS.n60 8.28285
R3833 VSS.n35 VSS.n14 8.28285
R3834 VSS.n956 VSS.t0 8.24205
R3835 VSS.n503 VSS.n498 8.2073
R3836 VSS.n442 VSS.n437 8.2073
R3837 VSS.n1642 VSS.n952 7.58273
R3838 VSS.n1640 VSS.n956 7.58273
R3839 VSS.n1649 VSS.n1648 7.58273
R3840 VSS.n1658 VSS.n1657 7.58273
R3841 VSS.n1666 VSS.n931 7.58273
R3842 VSS.n1664 VSS.n935 7.58273
R3843 VSS.n1674 VSS.t127 7.58273
R3844 VSS.n1673 VSS.n1672 7.58273
R3845 VSS.n1682 VSS.n1681 7.58273
R3846 VSS.n1690 VSS.n910 7.58273
R3847 VSS.n2053 VSS.n735 7.58273
R3848 VSS.n2006 VSS.n2005 7.52991
R3849 VSS.n1698 VSS.t4 7.25307
R3850 VSS.n838 VSS.t9 7.25307
R3851 VSS.n1531 VSS.t38 6.9234
R3852 VSS.t62 VSS.n918 6.9234
R3853 VSS.n176 VSS.n159 6.77697
R3854 VSS.n133 VSS.n132 6.77697
R3855 VSS.n76 VSS.n75 6.77697
R3856 VSS.n34 VSS.n16 6.77697
R3857 VSS.n1634 VSS.n960 6.59374
R3858 VSS.n1688 VSS.t1 6.59374
R3859 VSS.n2137 VSS.t128 6.59374
R3860 VSS.t98 VSS.n579 6.59374
R3861 VSS.n522 VSS.n509 6.41949
R3862 VSS.n519 VSS.n518 6.41949
R3863 VSS.n460 VSS.n459 6.41949
R3864 VSS.n462 VSS.n449 6.41949
R3865 VSS.n705 VSS.n702 6.41949
R3866 VSS.n678 VSS.n659 6.41949
R3867 VSS.n2369 VSS.n305 6.32304
R3868 VSS.n1501 VSS.t68 6.26408
R3869 VSS.t22 VSS.n791 6.26408
R3870 VSS.n2390 VSS.n100 6.14552
R3871 VSS.n2313 VSS.n2312 5.93442
R3872 VSS.n2003 VSS.n838 5.93442
R3873 VSS.n2306 VSS.n340 5.93442
R3874 VSS.n2251 VSS.n343 5.93442
R3875 VSS.n2389 VSS.n200 5.868
R3876 VSS.n526 VSS.t77 5.8005
R3877 VSS.n526 VSS.t32 5.8005
R3878 VSS.n517 VSS.t111 5.8005
R3879 VSS.n517 VSS.t77 5.8005
R3880 VSS.n504 VSS.t112 5.8005
R3881 VSS.n504 VSS.t13 5.8005
R3882 VSS.n452 VSS.t52 5.8005
R3883 VSS.n452 VSS.t50 5.8005
R3884 VSS.n466 VSS.t50 5.8005
R3885 VSS.n466 VSS.t110 5.8005
R3886 VSS.n443 VSS.t36 5.8005
R3887 VSS.n443 VSS.t94 5.8005
R3888 VSS.n490 VSS.t118 5.8005
R3889 VSS.n490 VSS.t107 5.8005
R3890 VSS.n486 VSS.t93 5.8005
R3891 VSS.n486 VSS.t109 5.8005
R3892 VSS.n482 VSS.t87 5.8005
R3893 VSS.n482 VSS.t96 5.8005
R3894 VSS.n478 VSS.t113 5.8005
R3895 VSS.n478 VSS.t83 5.8005
R3896 VSS.n474 VSS.t117 5.8005
R3897 VSS.n474 VSS.t115 5.8005
R3898 VSS.n470 VSS.t104 5.8005
R3899 VSS.n470 VSS.t92 5.8005
R3900 VSS.n488 VSS.t114 5.8005
R3901 VSS.n488 VSS.t84 5.8005
R3902 VSS.n484 VSS.t101 5.8005
R3903 VSS.n484 VSS.t100 5.8005
R3904 VSS.n480 VSS.t90 5.8005
R3905 VSS.n480 VSS.t91 5.8005
R3906 VSS.n476 VSS.t122 5.8005
R3907 VSS.n476 VSS.t121 5.8005
R3908 VSS.n472 VSS.t99 5.8005
R3909 VSS.n472 VSS.t82 5.8005
R3910 VSS.n711 VSS.t119 5.8005
R3911 VSS.t10 VSS.n711 5.8005
R3912 VSS.n712 VSS.t10 5.8005
R3913 VSS.n712 VSS.t44 5.8005
R3914 VSS.n694 VSS.t120 5.8005
R3915 VSS.n694 VSS.t89 5.8005
R3916 VSS.n692 VSS.t108 5.8005
R3917 VSS.n692 VSS.t102 5.8005
R3918 VSS.n690 VSS.t95 5.8005
R3919 VSS.n690 VSS.t97 5.8005
R3920 VSS.n688 VSS.t86 5.8005
R3921 VSS.n688 VSS.t85 5.8005
R3922 VSS.n686 VSS.t105 5.8005
R3923 VSS.n686 VSS.t88 5.8005
R3924 VSS.n682 VSS.t58 5.8005
R3925 VSS.n682 VSS.t116 5.8005
R3926 VSS.n675 VSS.t60 5.8005
R3927 VSS.n675 VSS.t58 5.8005
R3928 VSS.n1781 VSS.n1780 5.60476
R3929 VSS.n1780 VSS.n806 5.60476
R3930 VSS.n2031 VSS.n809 5.60476
R3931 VSS.n1801 VSS.n1800 5.60476
R3932 VSS.n1800 VSS.n1799 5.60476
R3933 VSS.n2025 VSS.n815 5.60476
R3934 VSS.n2025 VSS.n2024 5.60476
R3935 VSS.n1992 VSS.n818 5.60476
R3936 VSS.n2018 VSS.n832 5.60476
R3937 VSS.n2018 VSS.t126 5.60476
R3938 VSS.n2017 VSS.n2012 5.60476
R3939 VSS.n2011 VSS.n332 5.60476
R3940 VSS.n2312 VSS.n334 5.60476
R3941 VSS.n2003 VSS.n2002 5.60476
R3942 VSS.n2306 VSS.n2305 5.60476
R3943 VSS.n2251 VSS.n2250 5.60476
R3944 VSS.n719 VSS.n715 5.37662
R3945 VSS.n674 VSS.n662 5.37662
R3946 VSS.n177 VSS.n157 5.27109
R3947 VSS.n129 VSS.n116 5.27109
R3948 VSS.n79 VSS.n58 5.27109
R3949 VSS.n31 VSS.n30 5.27109
R3950 VSS.n1414 VSS.t103 4.94543
R3951 VSS.n1491 VSS.t68 4.94543
R3952 VSS.n1788 VSS.t22 4.94543
R3953 VSS.n1991 VSS.t106 4.94543
R3954 VSS.n2391 VSS.n0 4.78621
R3955 VSS.n1634 VSS.n1568 4.61577
R3956 VSS.n431 VSS.n389 4.51815
R3957 VSS.n1476 VSS.t38 4.28611
R3958 VSS.n1672 VSS.t62 4.28611
R3959 VSS.n2058 VSS.n2057 4.03565
R3960 VSS.t2 VSS.n2031 3.95645
R3961 VSS.n685 VSS.n656 3.81995
R3962 VSS.n181 VSS.n180 3.76521
R3963 VSS.n128 VSS.n118 3.76521
R3964 VSS.n525 VSS.n508 3.76521
R3965 VSS.n515 VSS.n512 3.76521
R3966 VSS.n495 VSS.n494 3.76521
R3967 VSS.n457 VSS.n456 3.76521
R3968 VSS.n465 VSS.n448 3.76521
R3969 VSS.n434 VSS.n433 3.76521
R3970 VSS.n722 VSS.n698 3.76521
R3971 VSS.n709 VSS.n703 3.76521
R3972 VSS.n681 VSS.n658 3.76521
R3973 VSS.n668 VSS.n667 3.76521
R3974 VSS.n913 VSS.n729 3.76521
R3975 VSS.n80 VSS.n56 3.76521
R3976 VSS.n27 VSS.n18 3.76521
R3977 VSS.t49 VSS.n1036 3.62678
R3978 VSS.n1554 VSS.n952 3.62678
R3979 VSS.n1641 VSS.n1640 3.62678
R3980 VSS.n1650 VSS.n1649 3.62678
R3981 VSS.n1658 VSS.n939 3.62678
R3982 VSS.n1656 VSS.n931 3.62678
R3983 VSS.n1665 VSS.n1664 3.62678
R3984 VSS.n935 VSS.t127 3.62678
R3985 VSS.n1674 VSS.n1673 3.62678
R3986 VSS.n1682 VSS.n918 3.62678
R3987 VSS.n1680 VSS.n910 3.62678
R3988 VSS.n1689 VSS.n1688 3.62678
R3989 VSS.n1699 VSS.n1698 3.62678
R3990 VSS.n2053 VSS.n734 3.62678
R3991 VSS.t9 VSS.n334 3.62678
R3992 VSS.n1414 VSS.n1026 3.29712
R3993 VSS.n1992 VSS.n1991 3.29712
R3994 VSS.n727 VSS.n0 3.163
R3995 VSS.n164 VSS.n162 3.09986
R3996 VSS.n144 VSS.n111 3.09986
R3997 VSS.n66 VSS.n65 3.09986
R3998 VSS.n41 VSS.n10 3.09986
R3999 VSS.n1650 VSS.t0 2.96746
R4000 VSS.n513 VSS.n492 2.89851
R4001 VSS.n469 VSS.n468 2.89851
R4002 VSS.n469 VSS.n446 2.82558
R4003 VSS.n2390 VSS.n2389 2.77891
R4004 VSS.n704 VSS.n696 2.67025
R4005 VSS.n726 VSS.n725 2.67025
R4006 VSS.n685 VSS.n684 2.67025
R4007 VSS.n2039 VSS.n797 2.6378
R4008 VSS.t23 VSS.n193 2.48621
R4009 VSS.n193 VSS.t16 2.48621
R4010 VSS.t81 VSS.n194 2.48621
R4011 VSS.n194 VSS.t23 2.48621
R4012 VSS.t63 VSS.n195 2.48621
R4013 VSS.n195 VSS.t81 2.48621
R4014 VSS.t66 VSS.n196 2.48621
R4015 VSS.n196 VSS.t63 2.48621
R4016 VSS.n145 VSS.t71 2.48621
R4017 VSS.t69 VSS.n145 2.48621
R4018 VSS.n146 VSS.t69 2.48621
R4019 VSS.n146 VSS.t7 2.48621
R4020 VSS.n149 VSS.t7 2.48621
R4021 VSS.t39 VSS.n149 2.48621
R4022 VSS.n150 VSS.t39 2.48621
R4023 VSS.t30 VSS.n150 2.48621
R4024 VSS.n197 VSS.t30 2.48621
R4025 VSS.n197 VSS.t66 2.48621
R4026 VSS.t47 VSS.n93 2.48621
R4027 VSS.n93 VSS.t41 2.48621
R4028 VSS.t25 VSS.n94 2.48621
R4029 VSS.n94 VSS.t47 2.48621
R4030 VSS.t73 VSS.n95 2.48621
R4031 VSS.n95 VSS.t25 2.48621
R4032 VSS.t75 VSS.n96 2.48621
R4033 VSS.n96 VSS.t73 2.48621
R4034 VSS.n45 VSS.t20 2.48621
R4035 VSS.t79 VSS.n45 2.48621
R4036 VSS.n46 VSS.t79 2.48621
R4037 VSS.n46 VSS.t27 2.48621
R4038 VSS.n49 VSS.t27 2.48621
R4039 VSS.t56 VSS.n49 2.48621
R4040 VSS.n50 VSS.t56 2.48621
R4041 VSS.t54 VSS.n50 2.48621
R4042 VSS.n97 VSS.t54 2.48621
R4043 VSS.n97 VSS.t75 2.48621
R4044 VSS.n2060 VSS.n2059 2.44251
R4045 VSS.n2058 VSS.n728 2.44179
R4046 VSS.n532 VSS.n531 2.33344
R4047 VSS.t29 VSS.n962 2.30813
R4048 VSS.t65 VSS.n939 2.30813
R4049 VSS.n184 VSS.n155 2.25932
R4050 VSS.n125 VSS.n124 2.25932
R4051 VSS.n499 VSS.n496 2.25932
R4052 VSS.n438 VSS.n435 2.25932
R4053 VSS.n721 VSS.n700 2.25932
R4054 VSS.n671 VSS.n663 2.25932
R4055 VSS.n84 VSS.n83 2.25932
R4056 VSS.n26 VSS.n20 2.25932
R4057 VSS.n530 VSS.n529 2.25177
R4058 VSS.n2391 VSS.n2390 1.73042
R4059 VSS.n1424 VSS.t19 1.64881
R4060 VSS.n2032 VSS.t2 1.64881
R4061 VSS.n687 VSS.n685 1.1502
R4062 VSS.n689 VSS.n687 1.1502
R4063 VSS.n691 VSS.n689 1.1502
R4064 VSS.n693 VSS.n691 1.1502
R4065 VSS.n695 VSS.n693 1.1502
R4066 VSS.n696 VSS.n695 1.1502
R4067 VSS.n726 VSS.n696 1.1502
R4068 VSS.n727 VSS.n726 1.01732
R4069 VSS.n2059 VSS.n2058 1.01577
R4070 VSS.t1 VSS.n903 0.989486
R4071 VSS.n1801 VSS.t124 0.989486
R4072 VSS.n2002 VSS.t3 0.989486
R4073 VSS.n2299 VSS.t12 0.989486
R4074 VSS.n531 VSS.n0 0.861992
R4075 VSS.n531 VSS.n530 0.7864
R4076 VSS.n192 VSS.n187 0.779912
R4077 VSS.n192 VSS.n152 0.779912
R4078 VSS.n152 VSS.n151 0.779912
R4079 VSS.n151 VSS.n104 0.779912
R4080 VSS.n121 VSS.n109 0.779912
R4081 VSS.n147 VSS.n109 0.779912
R4082 VSS.n148 VSS.n147 0.779912
R4083 VSS.n148 VSS.n103 0.779912
R4084 VSS.n198 VSS.n103 0.779912
R4085 VSS.n198 VSS.n104 0.779912
R4086 VSS.n92 VSS.n87 0.779912
R4087 VSS.n92 VSS.n52 0.779912
R4088 VSS.n52 VSS.n51 0.779912
R4089 VSS.n51 VSS.n4 0.779912
R4090 VSS.n21 VSS.n9 0.779912
R4091 VSS.n47 VSS.n9 0.779912
R4092 VSS.n48 VSS.n47 0.779912
R4093 VSS.n48 VSS.n3 0.779912
R4094 VSS.n98 VSS.n3 0.779912
R4095 VSS.n98 VSS.n4 0.779912
R4096 VSS.n718 VSS.n717 0.753441
R4097 VSS.n673 VSS.n672 0.753441
R4098 VSS.n2056 VSS.n730 0.753441
R4099 VSS.n188 VSS.n101 0.701719
R4100 VSS.n189 VSS.n188 0.701719
R4101 VSS.n190 VSS.n189 0.701719
R4102 VSS.n107 VSS.n106 0.701719
R4103 VSS.n106 VSS.n105 0.701719
R4104 VSS.n105 VSS.n102 0.701719
R4105 VSS.n88 VSS.n1 0.701719
R4106 VSS.n89 VSS.n88 0.701719
R4107 VSS.n90 VSS.n89 0.701719
R4108 VSS.n7 VSS.n6 0.701719
R4109 VSS.n6 VSS.n5 0.701719
R4110 VSS.n5 VSS.n2 0.701719
R4111 VSS.n1049 VSS.t35 0.659824
R4112 VSS.n2046 VSS.n741 0.659824
R4113 VSS.n529 VSS.n528 0.647239
R4114 VSS.n454 VSS.n446 0.647239
R4115 VSS.n471 VSS.n469 0.574311
R4116 VSS.n473 VSS.n471 0.574311
R4117 VSS.n475 VSS.n473 0.574311
R4118 VSS.n477 VSS.n475 0.574311
R4119 VSS.n479 VSS.n477 0.574311
R4120 VSS.n481 VSS.n479 0.574311
R4121 VSS.n483 VSS.n481 0.574311
R4122 VSS.n485 VSS.n483 0.574311
R4123 VSS.n487 VSS.n485 0.574311
R4124 VSS.n489 VSS.n487 0.574311
R4125 VSS.n491 VSS.n489 0.574311
R4126 VSS.n492 VSS.n491 0.574311
R4127 VSS.n530 VSS.n492 0.574311
R4128 VSS VSS.n2391 0.469656
R4129 VSS.n529 VSS.n506 0.418978
R4130 VSS.n446 VSS.n445 0.418978
R4131 VSS.n191 VSS.n190 0.35111
R4132 VSS.n108 VSS.n107 0.35111
R4133 VSS.n91 VSS.n90 0.35111
R4134 VSS.n8 VSS.n7 0.35111
R4135 VSS.n1050 VSS.n1049 0.330162
R4136 VSS.n1517 VSS.t6 0.330162
R4137 VSS.t4 VSS.n1697 0.330162
R4138 VSS.n2059 VSS.n727 0.32859
R4139 VSS.n520 VSS.n519 0.320353
R4140 VSS.n522 VSS.n520 0.320353
R4141 VSS.n522 VSS.n521 0.320353
R4142 VSS.n498 VSS.n497 0.320353
R4143 VSS.n462 VSS.n461 0.320353
R4144 VSS.n460 VSS.n450 0.320353
R4145 VSS.n461 VSS.n460 0.320353
R4146 VSS.n437 VSS.n436 0.320353
R4147 VSS.n705 VSS.n701 0.320353
R4148 VSS.n713 VSS.n701 0.320353
R4149 VSS.n714 VSS.n713 0.320353
R4150 VSS.n719 VSS.n714 0.320353
R4151 VSS.n662 VSS.n660 0.320353
R4152 VSS.n676 VSS.n660 0.320353
R4153 VSS.n677 VSS.n676 0.320353
R4154 VSS.n678 VSS.n677 0.320353
R4155 VSS.n199 VSS.n198 0.272321
R4156 VSS.n99 VSS.n98 0.272321
R4157 VSS.n199 VSS.n101 0.261436
R4158 VSS.n199 VSS.n102 0.261436
R4159 VSS.n99 VSS.n1 0.261436
R4160 VSS.n99 VSS.n2 0.261436
R4161 VSS.n192 VSS.n191 0.228761
R4162 VSS.n109 VSS.n108 0.228761
R4163 VSS.n92 VSS.n91 0.228761
R4164 VSS.n9 VSS.n8 0.228761
R4165 VSS.n187 VSS.n186 0.196152
R4166 VSS.n186 VSS.n154 0.196152
R4167 VSS.n179 VSS.n154 0.196152
R4168 VSS.n179 VSS.n178 0.196152
R4169 VSS.n178 VSS.n158 0.196152
R4170 VSS.n171 VSS.n158 0.196152
R4171 VSS.n171 VSS.n170 0.196152
R4172 VSS.n170 VSS.n162 0.196152
R4173 VSS.n121 VSS.n119 0.196152
R4174 VSS.n126 VSS.n119 0.196152
R4175 VSS.n127 VSS.n126 0.196152
R4176 VSS.n127 VSS.n115 0.196152
R4177 VSS.n134 VSS.n115 0.196152
R4178 VSS.n136 VSS.n134 0.196152
R4179 VSS.n136 VSS.n135 0.196152
R4180 VSS.n135 VSS.n111 0.196152
R4181 VSS.n514 VSS.n513 0.196152
R4182 VSS.n514 VSS.n510 0.196152
R4183 VSS.n519 VSS.n510 0.196152
R4184 VSS.n501 VSS.n498 0.196152
R4185 VSS.n501 VSS.n500 0.196152
R4186 VSS.n500 VSS.n493 0.196152
R4187 VSS.n506 VSS.n493 0.196152
R4188 VSS.n528 VSS.n507 0.196152
R4189 VSS.n523 VSS.n507 0.196152
R4190 VSS.n523 VSS.n522 0.196152
R4191 VSS.n468 VSS.n447 0.196152
R4192 VSS.n463 VSS.n447 0.196152
R4193 VSS.n463 VSS.n462 0.196152
R4194 VSS.n440 VSS.n437 0.196152
R4195 VSS.n440 VSS.n439 0.196152
R4196 VSS.n439 VSS.n432 0.196152
R4197 VSS.n445 VSS.n432 0.196152
R4198 VSS.n455 VSS.n454 0.196152
R4199 VSS.n455 VSS.n451 0.196152
R4200 VSS.n460 VSS.n451 0.196152
R4201 VSS.n708 VSS.n704 0.196152
R4202 VSS.n708 VSS.n707 0.196152
R4203 VSS.n707 VSS.n705 0.196152
R4204 VSS.n725 VSS.n697 0.196152
R4205 VSS.n720 VSS.n697 0.196152
R4206 VSS.n720 VSS.n719 0.196152
R4207 VSS.n666 VSS.n656 0.196152
R4208 VSS.n666 VSS.n665 0.196152
R4209 VSS.n665 VSS.n662 0.196152
R4210 VSS.n684 VSS.n657 0.196152
R4211 VSS.n679 VSS.n657 0.196152
R4212 VSS.n679 VSS.n678 0.196152
R4213 VSS.n66 VSS.n61 0.196152
R4214 VSS.n73 VSS.n61 0.196152
R4215 VSS.n74 VSS.n73 0.196152
R4216 VSS.n74 VSS.n57 0.196152
R4217 VSS.n81 VSS.n57 0.196152
R4218 VSS.n82 VSS.n81 0.196152
R4219 VSS.n82 VSS.n53 0.196152
R4220 VSS.n87 VSS.n53 0.196152
R4221 VSS.n41 VSS.n40 0.196152
R4222 VSS.n40 VSS.n13 0.196152
R4223 VSS.n33 VSS.n13 0.196152
R4224 VSS.n33 VSS.n32 0.196152
R4225 VSS.n32 VSS.n17 0.196152
R4226 VSS.n25 VSS.n17 0.196152
R4227 VSS.n25 VSS.n24 0.196152
R4228 VSS.n24 VSS.n21 0.196152
R4229 VSS.n200 VSS.n199 0.114136
R4230 VSS.n100 VSS.n99 0.114136
R4231 a_6681_4767.n49 a_6681_4767.n48 185
R4232 a_6681_4767.n48 a_6681_4767.n47 185
R4233 a_6681_4767.n48 a_6681_4767.n8 185
R4234 a_6681_4767.n48 a_6681_4767.n7 185
R4235 a_6681_4767.n48 a_6681_4767.n6 185
R4236 a_6681_4767.n48 a_6681_4767.n5 185
R4237 a_6681_4767.n48 a_6681_4767.n4 185
R4238 a_6681_4767.t2 a_6681_4767.n54 180.167
R4239 a_6681_4767.t2 a_6681_4767.n54 180.167
R4240 a_6681_4767.n53 a_6681_4767.t0 130.75
R4241 a_6681_4767.n48 a_6681_4767.n3 86.5152
R4242 a_6681_4767.n50 a_6681_4767.n0 30.3012
R4243 a_6681_4767.n31 a_6681_4767.n12 25.7063
R4244 a_6681_4767.n32 a_6681_4767.n11 25.7063
R4245 a_6681_4767.n10 a_6681_4767.n9 25.7063
R4246 a_6681_4767.n22 a_6681_4767.n21 25.7063
R4247 a_6681_4767.n23 a_6681_4767.n20 25.7063
R4248 a_6681_4767.n24 a_6681_4767.n19 25.7063
R4249 a_6681_4767.n25 a_6681_4767.n18 25.4781
R4250 a_6681_4767.n26 a_6681_4767.n17 25.4781
R4251 a_6681_4767.n27 a_6681_4767.n16 25.4781
R4252 a_6681_4767.n28 a_6681_4767.n15 25.4781
R4253 a_6681_4767.n29 a_6681_4767.n14 25.4781
R4254 a_6681_4767.n30 a_6681_4767.n13 25.4781
R4255 a_6681_4767.n35 a_6681_4767.n4 24.8476
R4256 a_6681_4767.n37 a_6681_4767.n5 23.3417
R4257 a_6681_4767.n34 a_6681_4767.n3 22.0256
R4258 a_6681_4767.n39 a_6681_4767.n6 21.8358
R4259 a_6681_4767.n41 a_6681_4767.n7 20.3299
R4260 a_6681_4767.n43 a_6681_4767.n8 18.824
R4261 a_6681_4767.n47 a_6681_4767.n46 17.3181
R4262 a_6681_4767.n48 a_6681_4767.n0 16.3559
R4263 a_6681_4767.n49 a_6681_4767.n2 15.8123
R4264 a_6681_4767.n35 a_6681_4767.n3 12.7256
R4265 a_6681_4767.n31 a_6681_4767.n30 12.3836
R4266 a_6681_4767.n25 a_6681_4767.n24 11.9167
R4267 a_6681_4767.n50 a_6681_4767.n49 11.2946
R4268 a_6681_4767.n47 a_6681_4767.n2 9.78874
R4269 a_6681_4767.n36 a_6681_4767.n35 9.3005
R4270 a_6681_4767.n38 a_6681_4767.n37 9.3005
R4271 a_6681_4767.n40 a_6681_4767.n39 9.3005
R4272 a_6681_4767.n42 a_6681_4767.n41 9.3005
R4273 a_6681_4767.n44 a_6681_4767.n43 9.3005
R4274 a_6681_4767.n46 a_6681_4767.n45 9.3005
R4275 a_6681_4767.n2 a_6681_4767.n1 9.3005
R4276 a_6681_4767.n51 a_6681_4767.n50 9.3005
R4277 a_6681_4767.n46 a_6681_4767.n8 8.28285
R4278 a_6681_4767.n43 a_6681_4767.n7 6.77697
R4279 a_6681_4767.n12 a_6681_4767.t8 5.8005
R4280 a_6681_4767.n12 a_6681_4767.t23 5.8005
R4281 a_6681_4767.n11 a_6681_4767.t17 5.8005
R4282 a_6681_4767.n11 a_6681_4767.t24 5.8005
R4283 a_6681_4767.n9 a_6681_4767.t12 5.8005
R4284 a_6681_4767.n9 a_6681_4767.t18 5.8005
R4285 a_6681_4767.n21 a_6681_4767.t5 5.8005
R4286 a_6681_4767.n21 a_6681_4767.t11 5.8005
R4287 a_6681_4767.n20 a_6681_4767.t7 5.8005
R4288 a_6681_4767.n20 a_6681_4767.t6 5.8005
R4289 a_6681_4767.n19 a_6681_4767.t22 5.8005
R4290 a_6681_4767.n19 a_6681_4767.t16 5.8005
R4291 a_6681_4767.n18 a_6681_4767.t19 5.8005
R4292 a_6681_4767.n18 a_6681_4767.t13 5.8005
R4293 a_6681_4767.n17 a_6681_4767.t3 5.8005
R4294 a_6681_4767.n17 a_6681_4767.t26 5.8005
R4295 a_6681_4767.n16 a_6681_4767.t25 5.8005
R4296 a_6681_4767.n16 a_6681_4767.t9 5.8005
R4297 a_6681_4767.n15 a_6681_4767.t10 5.8005
R4298 a_6681_4767.n15 a_6681_4767.t15 5.8005
R4299 a_6681_4767.n14 a_6681_4767.t14 5.8005
R4300 a_6681_4767.n14 a_6681_4767.t21 5.8005
R4301 a_6681_4767.n13 a_6681_4767.t4 5.8005
R4302 a_6681_4767.n13 a_6681_4767.t20 5.8005
R4303 a_6681_4767.n41 a_6681_4767.n6 5.27109
R4304 a_6681_4767.n39 a_6681_4767.n5 3.76521
R4305 a_6681_4767.n48 a_6681_4767.t27 2.48621
R4306 a_6681_4767.n48 a_6681_4767.t1 2.48621
R4307 a_6681_4767.n52 a_6681_4767.n0 2.36936
R4308 a_6681_4767.n37 a_6681_4767.n4 2.25932
R4309 a_6681_4767.n54 a_6681_4767.n53 1.27148
R4310 a_6681_4767.n26 a_6681_4767.n25 1.15229
R4311 a_6681_4767.n27 a_6681_4767.n26 1.15229
R4312 a_6681_4767.n28 a_6681_4767.n27 1.15229
R4313 a_6681_4767.n29 a_6681_4767.n28 1.15229
R4314 a_6681_4767.n30 a_6681_4767.n29 1.15229
R4315 a_6681_4767.n24 a_6681_4767.n23 1.15229
R4316 a_6681_4767.n23 a_6681_4767.n22 1.15229
R4317 a_6681_4767.n22 a_6681_4767.n10 1.15229
R4318 a_6681_4767.n32 a_6681_4767.n31 1.15229
R4319 a_6681_4767.n34 a_6681_4767.n33 0.791261
R4320 a_6681_4767.n33 a_6681_4767.n32 0.732643
R4321 a_6681_4767.n33 a_6681_4767.n10 0.420143
R4322 a_6681_4767.n53 a_6681_4767.n52 0.320353
R4323 a_6681_4767.n52 a_6681_4767.n51 0.196152
R4324 a_6681_4767.n51 a_6681_4767.n1 0.196152
R4325 a_6681_4767.n45 a_6681_4767.n1 0.196152
R4326 a_6681_4767.n45 a_6681_4767.n44 0.196152
R4327 a_6681_4767.n44 a_6681_4767.n42 0.196152
R4328 a_6681_4767.n42 a_6681_4767.n40 0.196152
R4329 a_6681_4767.n40 a_6681_4767.n38 0.196152
R4330 a_6681_4767.n38 a_6681_4767.n36 0.196152
R4331 a_6681_4767.n36 a_6681_4767.n34 0.196152
R4332 a_6681_14134.n69 a_6681_14134.t11 260.111
R4333 a_6681_14134.n67 a_6681_14134.t9 260.111
R4334 a_6681_14134.n70 a_6681_14134.t23 260.111
R4335 a_6681_14134.n65 a_6681_14134.t22 260.111
R4336 a_6681_14134.n67 a_6681_14134.t24 260.111
R4337 a_6681_14134.n69 a_6681_14134.t21 260.111
R4338 a_6681_14134.n70 a_6681_14134.t2 260.111
R4339 a_6681_14134.n65 a_6681_14134.t0 260.111
R4340 a_6681_14134.n68 a_6681_14134.n66 203.413
R4341 a_6681_14134.n72 a_6681_14134.n71 203.412
R4342 a_6681_14134.n29 a_6681_14134.n28 185
R4343 a_6681_14134.n29 a_6681_14134.n11 185
R4344 a_6681_14134.n29 a_6681_14134.n10 185
R4345 a_6681_14134.n29 a_6681_14134.n9 185
R4346 a_6681_14134.n29 a_6681_14134.n8 185
R4347 a_6681_14134.n29 a_6681_14134.n7 185
R4348 a_6681_14134.n29 a_6681_14134.n6 185
R4349 a_6681_14134.n60 a_6681_14134.n59 185
R4350 a_6681_14134.n60 a_6681_14134.n42 185
R4351 a_6681_14134.n60 a_6681_14134.n41 185
R4352 a_6681_14134.n60 a_6681_14134.n40 185
R4353 a_6681_14134.n60 a_6681_14134.n39 185
R4354 a_6681_14134.n60 a_6681_14134.n38 185
R4355 a_6681_14134.n60 a_6681_14134.n37 185
R4356 a_6681_14134.n12 a_6681_14134.t4 130.75
R4357 a_6681_14134.n43 a_6681_14134.t7 130.75
R4358 a_6681_14134.n12 a_6681_14134.t6 91.3557
R4359 a_6681_14134.n43 a_6681_14134.t8 91.3557
R4360 a_6681_14134.n30 a_6681_14134.n29 86.5152
R4361 a_6681_14134.n61 a_6681_14134.n60 86.5152
R4362 a_6681_14134.n14 a_6681_14134.n5 30.3012
R4363 a_6681_14134.n45 a_6681_14134.n36 30.3012
R4364 a_6681_14134.n66 a_6681_14134.t12 28.5655
R4365 a_6681_14134.n66 a_6681_14134.t10 28.5655
R4366 a_6681_14134.t1 a_6681_14134.n72 28.5655
R4367 a_6681_14134.n72 a_6681_14134.t3 28.5655
R4368 a_6681_14134.n28 a_6681_14134.n4 24.8476
R4369 a_6681_14134.n59 a_6681_14134.n35 24.8476
R4370 a_6681_14134.n27 a_6681_14134.n11 23.3417
R4371 a_6681_14134.n58 a_6681_14134.n42 23.3417
R4372 a_6681_14134.n31 a_6681_14134.n30 22.0256
R4373 a_6681_14134.n62 a_6681_14134.n61 22.0256
R4374 a_6681_14134.n24 a_6681_14134.n10 21.8358
R4375 a_6681_14134.n55 a_6681_14134.n41 21.8358
R4376 a_6681_14134.n22 a_6681_14134.n9 20.3299
R4377 a_6681_14134.n53 a_6681_14134.n40 20.3299
R4378 a_6681_14134.n20 a_6681_14134.n8 18.824
R4379 a_6681_14134.n51 a_6681_14134.n39 18.824
R4380 a_6681_14134.n2 a_6681_14134.n0 17.4823
R4381 a_6681_14134.n18 a_6681_14134.n7 17.3181
R4382 a_6681_14134.n49 a_6681_14134.n38 17.3181
R4383 a_6681_14134.n29 a_6681_14134.n5 16.3559
R4384 a_6681_14134.n60 a_6681_14134.n36 16.3559
R4385 a_6681_14134.n16 a_6681_14134.n6 15.8123
R4386 a_6681_14134.n47 a_6681_14134.n37 15.8123
R4387 a_6681_14134.n2 a_6681_14134.n1 14.6053
R4388 a_6681_14134.n33 a_6681_14134.n32 14.377
R4389 a_6681_14134.n30 a_6681_14134.n4 12.7256
R4390 a_6681_14134.n61 a_6681_14134.n35 12.7256
R4391 a_6681_14134.n65 a_6681_14134.n64 12.1798
R4392 a_6681_14134.n14 a_6681_14134.n6 11.2946
R4393 a_6681_14134.n45 a_6681_14134.n37 11.2946
R4394 a_6681_14134.n64 a_6681_14134.n2 10.4849
R4395 a_6681_14134.n16 a_6681_14134.n7 9.78874
R4396 a_6681_14134.n47 a_6681_14134.n38 9.78874
R4397 a_6681_14134.n4 a_6681_14134.n3 9.3005
R4398 a_6681_14134.n27 a_6681_14134.n26 9.3005
R4399 a_6681_14134.n25 a_6681_14134.n24 9.3005
R4400 a_6681_14134.n23 a_6681_14134.n22 9.3005
R4401 a_6681_14134.n21 a_6681_14134.n20 9.3005
R4402 a_6681_14134.n19 a_6681_14134.n18 9.3005
R4403 a_6681_14134.n17 a_6681_14134.n16 9.3005
R4404 a_6681_14134.n15 a_6681_14134.n14 9.3005
R4405 a_6681_14134.n35 a_6681_14134.n34 9.3005
R4406 a_6681_14134.n58 a_6681_14134.n57 9.3005
R4407 a_6681_14134.n56 a_6681_14134.n55 9.3005
R4408 a_6681_14134.n54 a_6681_14134.n53 9.3005
R4409 a_6681_14134.n52 a_6681_14134.n51 9.3005
R4410 a_6681_14134.n50 a_6681_14134.n49 9.3005
R4411 a_6681_14134.n48 a_6681_14134.n47 9.3005
R4412 a_6681_14134.n46 a_6681_14134.n45 9.3005
R4413 a_6681_14134.n18 a_6681_14134.n8 8.28285
R4414 a_6681_14134.n49 a_6681_14134.n39 8.28285
R4415 a_6681_14134.n20 a_6681_14134.n9 6.77697
R4416 a_6681_14134.n51 a_6681_14134.n40 6.77697
R4417 a_6681_14134.n33 a_6681_14134.n31 6.19091
R4418 a_6681_14134.n22 a_6681_14134.n10 5.27109
R4419 a_6681_14134.n53 a_6681_14134.n41 5.27109
R4420 a_6681_14134.n24 a_6681_14134.n11 3.76521
R4421 a_6681_14134.n55 a_6681_14134.n42 3.76521
R4422 a_6681_14134.n63 a_6681_14134.n62 3.31388
R4423 a_6681_14134.n0 a_6681_14134.t13 2.48621
R4424 a_6681_14134.n0 a_6681_14134.t15 2.48621
R4425 a_6681_14134.n1 a_6681_14134.t18 2.48621
R4426 a_6681_14134.n1 a_6681_14134.t16 2.48621
R4427 a_6681_14134.n29 a_6681_14134.t19 2.48621
R4428 a_6681_14134.n29 a_6681_14134.t5 2.48621
R4429 a_6681_14134.n32 a_6681_14134.t17 2.48621
R4430 a_6681_14134.n32 a_6681_14134.t14 2.48621
R4431 a_6681_14134.n60 a_6681_14134.t8 2.48621
R4432 a_6681_14134.n60 a_6681_14134.t20 2.48621
R4433 a_6681_14134.n13 a_6681_14134.n5 2.36936
R4434 a_6681_14134.n44 a_6681_14134.n36 2.36936
R4435 a_6681_14134.n63 a_6681_14134.n33 2.30287
R4436 a_6681_14134.n28 a_6681_14134.n27 2.25932
R4437 a_6681_14134.n59 a_6681_14134.n58 2.25932
R4438 a_6681_14134.n64 a_6681_14134.n63 1.07418
R4439 a_6681_14134.n13 a_6681_14134.n12 0.320353
R4440 a_6681_14134.n44 a_6681_14134.n43 0.320353
R4441 a_6681_14134.n31 a_6681_14134.n3 0.196152
R4442 a_6681_14134.n26 a_6681_14134.n3 0.196152
R4443 a_6681_14134.n26 a_6681_14134.n25 0.196152
R4444 a_6681_14134.n25 a_6681_14134.n23 0.196152
R4445 a_6681_14134.n23 a_6681_14134.n21 0.196152
R4446 a_6681_14134.n21 a_6681_14134.n19 0.196152
R4447 a_6681_14134.n19 a_6681_14134.n17 0.196152
R4448 a_6681_14134.n17 a_6681_14134.n15 0.196152
R4449 a_6681_14134.n15 a_6681_14134.n13 0.196152
R4450 a_6681_14134.n62 a_6681_14134.n34 0.196152
R4451 a_6681_14134.n57 a_6681_14134.n34 0.196152
R4452 a_6681_14134.n57 a_6681_14134.n56 0.196152
R4453 a_6681_14134.n56 a_6681_14134.n54 0.196152
R4454 a_6681_14134.n54 a_6681_14134.n52 0.196152
R4455 a_6681_14134.n52 a_6681_14134.n50 0.196152
R4456 a_6681_14134.n50 a_6681_14134.n48 0.196152
R4457 a_6681_14134.n48 a_6681_14134.n46 0.196152
R4458 a_6681_14134.n46 a_6681_14134.n44 0.196152
R4459 a_6681_14134.n70 a_6681_14134.n69 0.0850588
R4460 a_6681_14134.n71 a_6681_14134.n65 0.0427794
R4461 a_6681_14134.n71 a_6681_14134.n70 0.0427794
R4462 a_6681_14134.n69 a_6681_14134.n68 0.0427794
R4463 a_6681_14134.n68 a_6681_14134.n67 0.0427794
R4464 VDD.n213 VDD.n120 723.529
R4465 VDD.n135 VDD.n123 723.529
R4466 VDD.n268 VDD.n65 723.529
R4467 VDD.n82 VDD.n70 723.529
R4468 VDD.n190 VDD.n189 515.294
R4469 VDD.n202 VDD.n201 275.295
R4470 VDD.n278 VDD.n277 275.295
R4471 VDD.n310 VDD.t56 260.486
R4472 VDD.n333 VDD.t36 260.486
R4473 VDD.n16 VDD.t40 260.486
R4474 VDD.n40 VDD.t58 260.486
R4475 VDD.t63 VDD.n307 260.298
R4476 VDD.t48 VDD.n309 260.298
R4477 VDD.n314 VDD.t63 260.298
R4478 VDD.n330 VDD.t66 260.298
R4479 VDD.t66 VDD.n327 260.298
R4480 VDD.n334 VDD.t52 260.298
R4481 VDD.t42 VDD.n20 260.298
R4482 VDD.n18 VDD.t31 260.298
R4483 VDD.n21 VDD.t42 260.298
R4484 VDD.t38 VDD.n39 260.298
R4485 VDD.n37 VDD.t46 260.298
R4486 VDD.n33 VDD.t46 260.298
R4487 VDD.n2 VDD.t60 260.199
R4488 VDD.n350 VDD.t28 260.199
R4489 VDD.n313 VDD.t26 260.111
R4490 VDD.t26 VDD.n312 260.111
R4491 VDD.n310 VDD.t48 260.111
R4492 VDD.t52 VDD.n333 260.111
R4493 VDD.n332 VDD.t33 260.111
R4494 VDD.t33 VDD.n331 260.111
R4495 VDD.t50 VDD.n14 260.111
R4496 VDD.n19 VDD.t50 260.111
R4497 VDD.t31 VDD.n16 260.111
R4498 VDD.n40 VDD.t38 260.111
R4499 VDD.t54 VDD.n32 260.111
R4500 VDD.n38 VDD.t54 260.111
R4501 VDD.n137 VDD.n136 240
R4502 VDD.n208 VDD.n136 240
R4503 VDD.n206 VDD.n205 240
R4504 VDD.n198 VDD.n197 240
R4505 VDD.n194 VDD.n193 240
R4506 VDD.n186 VDD.n185 240
R4507 VDD.n182 VDD.n181 240
R4508 VDD.n178 VDD.n177 240
R4509 VDD.n174 VDD.n173 240
R4510 VDD.n170 VDD.n169 240
R4511 VDD.n166 VDD.n135 240
R4512 VDD.n264 VDD.n65 240
R4513 VDD.n264 VDD.n67 240
R4514 VDD.n87 VDD.n67 240
R4515 VDD.n88 VDD.n87 240
R4516 VDD.n89 VDD.n88 240
R4517 VDD.n141 VDD.n89 240
R4518 VDD.n141 VDD.n94 240
R4519 VDD.n95 VDD.n94 240
R4520 VDD.n96 VDD.n95 240
R4521 VDD.n146 VDD.n96 240
R4522 VDD.n146 VDD.n101 240
R4523 VDD.n102 VDD.n101 240
R4524 VDD.n103 VDD.n102 240
R4525 VDD.n151 VDD.n103 240
R4526 VDD.n151 VDD.n108 240
R4527 VDD.n109 VDD.n108 240
R4528 VDD.n110 VDD.n109 240
R4529 VDD.n156 VDD.n110 240
R4530 VDD.n156 VDD.n115 240
R4531 VDD.n116 VDD.n115 240
R4532 VDD.n117 VDD.n116 240
R4533 VDD.n161 VDD.n117 240
R4534 VDD.n161 VDD.n122 240
R4535 VDD.n123 VDD.n122 240
R4536 VDD.n80 VDD.n79 240
R4537 VDD.n77 VDD.n75 240
R4538 VDD.n301 VDD.n49 240
R4539 VDD.n299 VDD.n298 240
R4540 VDD.n296 VDD.n53 240
R4541 VDD.n292 VDD.n291 240
R4542 VDD.n289 VDD.n56 240
R4543 VDD.n285 VDD.n284 240
R4544 VDD.n282 VDD.n59 240
R4545 VDD.n275 VDD.n62 240
R4546 VDD.n271 VDD.n270 240
R4547 VDD.n262 VDD.n70 240
R4548 VDD.n262 VDD.n71 240
R4549 VDD.n258 VDD.n71 240
R4550 VDD.n258 VDD.n86 240
R4551 VDD.n254 VDD.n86 240
R4552 VDD.n254 VDD.n91 240
R4553 VDD.n250 VDD.n91 240
R4554 VDD.n250 VDD.n93 240
R4555 VDD.n246 VDD.n93 240
R4556 VDD.n246 VDD.n98 240
R4557 VDD.n242 VDD.n98 240
R4558 VDD.n242 VDD.n100 240
R4559 VDD.n238 VDD.n100 240
R4560 VDD.n238 VDD.n104 240
R4561 VDD.n234 VDD.n104 240
R4562 VDD.n234 VDD.n106 240
R4563 VDD.n230 VDD.n106 240
R4564 VDD.n230 VDD.n111 240
R4565 VDD.n226 VDD.n111 240
R4566 VDD.n226 VDD.n113 240
R4567 VDD.n222 VDD.n113 240
R4568 VDD.n222 VDD.n118 240
R4569 VDD.n218 VDD.n118 240
R4570 VDD.n218 VDD.n120 240
R4571 VDD.n315 VDD.t65 232.03
R4572 VDD.t67 VDD.n326 232.03
R4573 VDD.n13 VDD.t45 232.03
R4574 VDD.n36 VDD.t47 232.03
R4575 VDD.n1 VDD.t62 231.756
R4576 VDD.n344 VDD.n342 206.48
R4577 VDD.n344 VDD.n343 205.865
R4578 VDD.n346 VDD.n345 205.865
R4579 VDD.n348 VDD.n347 205.865
R4580 VDD.n323 VDD.n322 205.865
R4581 VDD.n4 VDD.n3 205.865
R4582 VDD.n6 VDD.n5 205.865
R4583 VDD.n8 VDD.n7 205.865
R4584 VDD.n10 VDD.n9 205.865
R4585 VDD.n29 VDD.n28 205.865
R4586 VDD.n1 VDD.n0 203.142
R4587 VDD.n321 VDD.n320 203.127
R4588 VDD.n340 VDD.n339 203.127
R4589 VDD.n27 VDD.n26 203.127
R4590 VDD.n46 VDD.n45 203.127
R4591 VDD.n319 VDD.n305 203.126
R4592 VDD.n338 VDD.n324 203.126
R4593 VDD.n25 VDD.n11 203.126
R4594 VDD.n44 VDD.n30 203.126
R4595 VDD.n318 VDD.n306 203.03
R4596 VDD.n317 VDD.n316 203.03
R4597 VDD.n337 VDD.n336 203.03
R4598 VDD.n329 VDD.n328 203.03
R4599 VDD.n24 VDD.n12 203.03
R4600 VDD.n23 VDD.n22 203.03
R4601 VDD.n43 VDD.n42 203.03
R4602 VDD.n35 VDD.n34 203.03
R4603 VDD.n84 VDD.n70 185
R4604 VDD.n70 VDD.n69 185
R4605 VDD.n262 VDD.n261 185
R4606 VDD.n263 VDD.n262 185
R4607 VDD.n260 VDD.n71 185
R4608 VDD.n71 VDD.n68 185
R4609 VDD.n259 VDD.n258 185
R4610 VDD.n258 VDD.n257 185
R4611 VDD.n86 VDD.n85 185
R4612 VDD.n256 VDD.n86 185
R4613 VDD.n254 VDD.n253 185
R4614 VDD.n255 VDD.n254 185
R4615 VDD.n252 VDD.n91 185
R4616 VDD.n91 VDD.n90 185
R4617 VDD.n251 VDD.n250 185
R4618 VDD.n250 VDD.n249 185
R4619 VDD.n93 VDD.n92 185
R4620 VDD.n248 VDD.n93 185
R4621 VDD.n246 VDD.n245 185
R4622 VDD.n247 VDD.n246 185
R4623 VDD.n244 VDD.n98 185
R4624 VDD.n98 VDD.n97 185
R4625 VDD.n243 VDD.n242 185
R4626 VDD.n242 VDD.n241 185
R4627 VDD.n100 VDD.n99 185
R4628 VDD.n240 VDD.n100 185
R4629 VDD.n238 VDD.n237 185
R4630 VDD.n239 VDD.n238 185
R4631 VDD.n236 VDD.n104 185
R4632 VDD.n107 VDD.n104 185
R4633 VDD.n235 VDD.n234 185
R4634 VDD.n234 VDD.n233 185
R4635 VDD.n106 VDD.n105 185
R4636 VDD.n232 VDD.n106 185
R4637 VDD.n230 VDD.n229 185
R4638 VDD.n231 VDD.n230 185
R4639 VDD.n228 VDD.n111 185
R4640 VDD.n114 VDD.n111 185
R4641 VDD.n227 VDD.n226 185
R4642 VDD.n226 VDD.n225 185
R4643 VDD.n113 VDD.n112 185
R4644 VDD.n224 VDD.n113 185
R4645 VDD.n222 VDD.n221 185
R4646 VDD.n223 VDD.n222 185
R4647 VDD.n220 VDD.n118 185
R4648 VDD.n121 VDD.n118 185
R4649 VDD.n219 VDD.n218 185
R4650 VDD.n218 VDD.n217 185
R4651 VDD.n120 VDD.n119 185
R4652 VDD.n216 VDD.n120 185
R4653 VDD.n213 VDD.n212 185
R4654 VDD.n211 VDD.n137 185
R4655 VDD.n210 VDD.n136 185
R4656 VDD.n215 VDD.n136 185
R4657 VDD.n209 VDD.n208 185
R4658 VDD.n207 VDD.n206 185
R4659 VDD.n205 VDD.n204 185
R4660 VDD.n203 VDD.n202 185
R4661 VDD.n201 VDD.n200 185
R4662 VDD.n199 VDD.n198 185
R4663 VDD.n197 VDD.n196 185
R4664 VDD.n195 VDD.n194 185
R4665 VDD.n193 VDD.n192 185
R4666 VDD.n191 VDD.n190 185
R4667 VDD.n189 VDD.n188 185
R4668 VDD.n187 VDD.n186 185
R4669 VDD.n185 VDD.n184 185
R4670 VDD.n183 VDD.n182 185
R4671 VDD.n181 VDD.n180 185
R4672 VDD.n179 VDD.n178 185
R4673 VDD.n177 VDD.n176 185
R4674 VDD.n175 VDD.n174 185
R4675 VDD.n173 VDD.n172 185
R4676 VDD.n171 VDD.n170 185
R4677 VDD.n169 VDD.n168 185
R4678 VDD.n167 VDD.n166 185
R4679 VDD.n165 VDD.n135 185
R4680 VDD.n215 VDD.n135 185
R4681 VDD.n164 VDD.n123 185
R4682 VDD.n216 VDD.n123 185
R4683 VDD.n163 VDD.n122 185
R4684 VDD.n217 VDD.n122 185
R4685 VDD.n162 VDD.n161 185
R4686 VDD.n161 VDD.n121 185
R4687 VDD.n160 VDD.n117 185
R4688 VDD.n223 VDD.n117 185
R4689 VDD.n159 VDD.n116 185
R4690 VDD.n224 VDD.n116 185
R4691 VDD.n158 VDD.n115 185
R4692 VDD.n225 VDD.n115 185
R4693 VDD.n157 VDD.n156 185
R4694 VDD.n156 VDD.n114 185
R4695 VDD.n155 VDD.n110 185
R4696 VDD.n231 VDD.n110 185
R4697 VDD.n154 VDD.n109 185
R4698 VDD.n232 VDD.n109 185
R4699 VDD.n153 VDD.n108 185
R4700 VDD.n233 VDD.n108 185
R4701 VDD.n152 VDD.n151 185
R4702 VDD.n151 VDD.n107 185
R4703 VDD.n150 VDD.n103 185
R4704 VDD.n239 VDD.n103 185
R4705 VDD.n149 VDD.n102 185
R4706 VDD.n240 VDD.n102 185
R4707 VDD.n148 VDD.n101 185
R4708 VDD.n241 VDD.n101 185
R4709 VDD.n147 VDD.n146 185
R4710 VDD.n146 VDD.n97 185
R4711 VDD.n145 VDD.n96 185
R4712 VDD.n247 VDD.n96 185
R4713 VDD.n144 VDD.n95 185
R4714 VDD.n248 VDD.n95 185
R4715 VDD.n143 VDD.n94 185
R4716 VDD.n249 VDD.n94 185
R4717 VDD.n142 VDD.n141 185
R4718 VDD.n141 VDD.n90 185
R4719 VDD.n140 VDD.n89 185
R4720 VDD.n255 VDD.n89 185
R4721 VDD.n139 VDD.n88 185
R4722 VDD.n256 VDD.n88 185
R4723 VDD.n138 VDD.n87 185
R4724 VDD.n257 VDD.n87 185
R4725 VDD.n67 VDD.n66 185
R4726 VDD.n68 VDD.n67 185
R4727 VDD.n265 VDD.n264 185
R4728 VDD.n264 VDD.n263 185
R4729 VDD.n266 VDD.n65 185
R4730 VDD.n69 VDD.n65 185
R4731 VDD.n268 VDD.n267 185
R4732 VDD.n270 VDD.n63 185
R4733 VDD.n272 VDD.n271 185
R4734 VDD.n273 VDD.n62 185
R4735 VDD.n275 VDD.n274 185
R4736 VDD.n277 VDD.n60 185
R4737 VDD.n279 VDD.n278 185
R4738 VDD.n280 VDD.n59 185
R4739 VDD.n282 VDD.n281 185
R4740 VDD.n284 VDD.n57 185
R4741 VDD.n286 VDD.n285 185
R4742 VDD.n287 VDD.n56 185
R4743 VDD.n289 VDD.n288 185
R4744 VDD.n291 VDD.n54 185
R4745 VDD.n293 VDD.n292 185
R4746 VDD.n294 VDD.n53 185
R4747 VDD.n296 VDD.n295 185
R4748 VDD.n298 VDD.n52 185
R4749 VDD.n299 VDD.n50 185
R4750 VDD.n302 VDD.n301 185
R4751 VDD.n303 VDD.n49 185
R4752 VDD.n75 VDD.n48 185
R4753 VDD.n77 VDD.n76 185
R4754 VDD.n79 VDD.n73 185
R4755 VDD.n80 VDD.n72 185
R4756 VDD.n83 VDD.n82 185
R4757 VDD.n290 VDD.n289 107.683
R4758 VDD.n291 VDD.n290 107.683
R4759 VDD.n350 VDD.n349 101.662
R4760 VDD.n177 VDD.n132 78.9253
R4761 VDD.n300 VDD.n299 78.9253
R4762 VDD.n174 VDD.n132 78.9253
R4763 VDD.n301 VDD.n300 78.9253
R4764 VDD.n84 VDD.n83 77.177
R4765 VDD.n212 VDD.n119 77.177
R4766 VDD.n165 VDD.n164 77.177
R4767 VDD.n267 VDD.n266 77.177
R4768 VDD.n214 VDD.n213 72.7879
R4769 VDD.n208 VDD.n124 72.7879
R4770 VDD.n205 VDD.n125 72.7879
R4771 VDD.n201 VDD.n126 72.7879
R4772 VDD.n197 VDD.n127 72.7879
R4773 VDD.n193 VDD.n128 72.7879
R4774 VDD.n189 VDD.n129 72.7879
R4775 VDD.n185 VDD.n130 72.7879
R4776 VDD.n181 VDD.n131 72.7879
R4777 VDD.n173 VDD.n133 72.7879
R4778 VDD.n169 VDD.n134 72.7879
R4779 VDD.n81 VDD.n80 72.7879
R4780 VDD.n78 VDD.n77 72.7879
R4781 VDD.n74 VDD.n49 72.7879
R4782 VDD.n297 VDD.n296 72.7879
R4783 VDD.n292 VDD.n55 72.7879
R4784 VDD.n285 VDD.n58 72.7879
R4785 VDD.n283 VDD.n282 72.7879
R4786 VDD.n278 VDD.n61 72.7879
R4787 VDD.n276 VDD.n275 72.7879
R4788 VDD.n271 VDD.n64 72.7879
R4789 VDD.n269 VDD.n268 72.7879
R4790 VDD.n214 VDD.n137 72.7879
R4791 VDD.n206 VDD.n124 72.7879
R4792 VDD.n202 VDD.n125 72.7879
R4793 VDD.n198 VDD.n126 72.7879
R4794 VDD.n194 VDD.n127 72.7879
R4795 VDD.n190 VDD.n128 72.7879
R4796 VDD.n186 VDD.n129 72.7879
R4797 VDD.n182 VDD.n130 72.7879
R4798 VDD.n178 VDD.n131 72.7879
R4799 VDD.n170 VDD.n133 72.7879
R4800 VDD.n166 VDD.n134 72.7879
R4801 VDD.n270 VDD.n269 72.7879
R4802 VDD.n64 VDD.n62 72.7879
R4803 VDD.n277 VDD.n276 72.7879
R4804 VDD.n61 VDD.n59 72.7879
R4805 VDD.n284 VDD.n283 72.7879
R4806 VDD.n58 VDD.n56 72.7879
R4807 VDD.n55 VDD.n53 72.7879
R4808 VDD.n298 VDD.n297 72.7879
R4809 VDD.n75 VDD.n74 72.7879
R4810 VDD.n79 VDD.n78 72.7879
R4811 VDD.n82 VDD.n81 72.7879
R4812 VDD.n69 VDD.n51 57.1093
R4813 VDD.n216 VDD.n215 57.1093
R4814 VDD.n215 VDD.n214 56.1076
R4815 VDD.n215 VDD.n124 56.1076
R4816 VDD.n215 VDD.n125 56.1076
R4817 VDD.n215 VDD.n126 56.1076
R4818 VDD.n215 VDD.n127 56.1076
R4819 VDD.n215 VDD.n128 56.1076
R4820 VDD.n215 VDD.n129 56.1076
R4821 VDD.n215 VDD.n130 56.1076
R4822 VDD.n215 VDD.n131 56.1076
R4823 VDD.n215 VDD.n133 56.1076
R4824 VDD.n215 VDD.n134 56.1076
R4825 VDD.n269 VDD.n51 56.1076
R4826 VDD.n64 VDD.n51 56.1076
R4827 VDD.n276 VDD.n51 56.1076
R4828 VDD.n61 VDD.n51 56.1076
R4829 VDD.n283 VDD.n51 56.1076
R4830 VDD.n58 VDD.n51 56.1076
R4831 VDD.n55 VDD.n51 56.1076
R4832 VDD.n297 VDD.n51 56.1076
R4833 VDD.n74 VDD.n51 56.1076
R4834 VDD.n78 VDD.n51 56.1076
R4835 VDD.n81 VDD.n51 56.1076
R4836 VDD.n191 VDD.n188 54.9652
R4837 VDD.n288 VDD.n54 54.9652
R4838 VDD.n215 VDD.n132 53.0388
R4839 VDD.n300 VDD.n51 53.0388
R4840 VDD.n349 VDD.t69 41.0864
R4841 VDD.n290 VDD.n51 38.6605
R4842 VDD.n263 VDD.n68 30.8211
R4843 VDD.n257 VDD.n256 30.8211
R4844 VDD.n255 VDD.n90 30.8211
R4845 VDD.n249 VDD.n248 30.8211
R4846 VDD.n247 VDD.n97 30.8211
R4847 VDD.n241 VDD.n240 30.8211
R4848 VDD.n240 VDD.n239 30.8211
R4849 VDD.n233 VDD.n107 30.8211
R4850 VDD.n232 VDD.n231 30.8211
R4851 VDD.n225 VDD.n114 30.8211
R4852 VDD.n224 VDD.n223 30.8211
R4853 VDD.n217 VDD.n121 30.8211
R4854 VDD.t0 VDD.n97 30.3679
R4855 VDD.n107 VDD.t14 30.3679
R4856 VDD.n248 VDD.t17 29.4614
R4857 VDD.t11 VDD.n232 29.4614
R4858 VDD.n203 VDD.n200 29.3652
R4859 VDD.n176 VDD.n175 29.3652
R4860 VDD.n302 VDD.n50 29.3652
R4861 VDD.n279 VDD.n60 29.3652
R4862 VDD.n0 VDD.t24 28.5655
R4863 VDD.n0 VDD.t61 28.5655
R4864 VDD.n3 VDD.t9 28.5655
R4865 VDD.n3 VDD.t10 28.5655
R4866 VDD.n5 VDD.t72 28.5655
R4867 VDD.n5 VDD.t71 28.5655
R4868 VDD.n7 VDD.t76 28.5655
R4869 VDD.n7 VDD.t1 28.5655
R4870 VDD.n9 VDD.t4 28.5655
R4871 VDD.n9 VDD.t23 28.5655
R4872 VDD.n342 VDD.t6 28.5655
R4873 VDD.n342 VDD.t8 28.5655
R4874 VDD.n343 VDD.t74 28.5655
R4875 VDD.n343 VDD.t25 28.5655
R4876 VDD.n345 VDD.t70 28.5655
R4877 VDD.n345 VDD.t75 28.5655
R4878 VDD.n347 VDD.t73 28.5655
R4879 VDD.n347 VDD.t68 28.5655
R4880 VDD.n320 VDD.t12 28.5655
R4881 VDD.n320 VDD.t57 28.5655
R4882 VDD.t49 VDD.n318 28.5655
R4883 VDD.n318 VDD.t27 28.5655
R4884 VDD.t27 VDD.n317 28.5655
R4885 VDD.n317 VDD.t64 28.5655
R4886 VDD.t57 VDD.n319 28.5655
R4887 VDD.n319 VDD.t49 28.5655
R4888 VDD.n339 VDD.t37 28.5655
R4889 VDD.n339 VDD.t21 28.5655
R4890 VDD.n337 VDD.t35 28.5655
R4891 VDD.t53 VDD.n337 28.5655
R4892 VDD.n328 VDD.t67 28.5655
R4893 VDD.n328 VDD.t35 28.5655
R4894 VDD.n338 VDD.t53 28.5655
R4895 VDD.t37 VDD.n338 28.5655
R4896 VDD.n322 VDD.t16 28.5655
R4897 VDD.n322 VDD.t19 28.5655
R4898 VDD.t32 VDD.n24 28.5655
R4899 VDD.n24 VDD.t51 28.5655
R4900 VDD.t51 VDD.n23 28.5655
R4901 VDD.n23 VDD.t44 28.5655
R4902 VDD.t41 VDD.n25 28.5655
R4903 VDD.n25 VDD.t32 28.5655
R4904 VDD.n26 VDD.t20 28.5655
R4905 VDD.n26 VDD.t41 28.5655
R4906 VDD.n28 VDD.t13 28.5655
R4907 VDD.n28 VDD.t15 28.5655
R4908 VDD.n43 VDD.t55 28.5655
R4909 VDD.t39 VDD.n43 28.5655
R4910 VDD.n34 VDD.t47 28.5655
R4911 VDD.n34 VDD.t55 28.5655
R4912 VDD.n44 VDD.t39 28.5655
R4913 VDD.t59 VDD.n44 28.5655
R4914 VDD.n45 VDD.t59 28.5655
R4915 VDD.n45 VDD.t18 28.5655
R4916 VDD.t22 VDD.n90 28.5549
R4917 VDD.n114 VDD.t5 28.5549
R4918 VDD.n256 VDD.t3 27.6484
R4919 VDD.t7 VDD.n224 27.6484
R4920 VDD.t34 VDD.n68 26.7419
R4921 VDD.n121 VDD.t2 26.7419
R4922 VDD.n69 VDD.t29 25.8354
R4923 VDD.t43 VDD.n216 25.8354
R4924 VDD.n261 VDD.n84 25.6005
R4925 VDD.n261 VDD.n260 25.6005
R4926 VDD.n260 VDD.n259 25.6005
R4927 VDD.n259 VDD.n85 25.6005
R4928 VDD.n253 VDD.n85 25.6005
R4929 VDD.n253 VDD.n252 25.6005
R4930 VDD.n252 VDD.n251 25.6005
R4931 VDD.n251 VDD.n92 25.6005
R4932 VDD.n245 VDD.n92 25.6005
R4933 VDD.n245 VDD.n244 25.6005
R4934 VDD.n244 VDD.n243 25.6005
R4935 VDD.n243 VDD.n99 25.6005
R4936 VDD.n237 VDD.n99 25.6005
R4937 VDD.n237 VDD.n236 25.6005
R4938 VDD.n236 VDD.n235 25.6005
R4939 VDD.n235 VDD.n105 25.6005
R4940 VDD.n229 VDD.n105 25.6005
R4941 VDD.n229 VDD.n228 25.6005
R4942 VDD.n228 VDD.n227 25.6005
R4943 VDD.n227 VDD.n112 25.6005
R4944 VDD.n221 VDD.n112 25.6005
R4945 VDD.n221 VDD.n220 25.6005
R4946 VDD.n220 VDD.n219 25.6005
R4947 VDD.n219 VDD.n119 25.6005
R4948 VDD.n212 VDD.n211 25.6005
R4949 VDD.n211 VDD.n210 25.6005
R4950 VDD.n210 VDD.n209 25.6005
R4951 VDD.n209 VDD.n207 25.6005
R4952 VDD.n207 VDD.n204 25.6005
R4953 VDD.n204 VDD.n203 25.6005
R4954 VDD.n200 VDD.n199 25.6005
R4955 VDD.n199 VDD.n196 25.6005
R4956 VDD.n196 VDD.n195 25.6005
R4957 VDD.n195 VDD.n192 25.6005
R4958 VDD.n192 VDD.n191 25.6005
R4959 VDD.n188 VDD.n187 25.6005
R4960 VDD.n187 VDD.n184 25.6005
R4961 VDD.n184 VDD.n183 25.6005
R4962 VDD.n183 VDD.n180 25.6005
R4963 VDD.n180 VDD.n179 25.6005
R4964 VDD.n179 VDD.n176 25.6005
R4965 VDD.n175 VDD.n172 25.6005
R4966 VDD.n172 VDD.n171 25.6005
R4967 VDD.n171 VDD.n168 25.6005
R4968 VDD.n168 VDD.n167 25.6005
R4969 VDD.n167 VDD.n165 25.6005
R4970 VDD.n266 VDD.n265 25.6005
R4971 VDD.n265 VDD.n66 25.6005
R4972 VDD.n138 VDD.n66 25.6005
R4973 VDD.n139 VDD.n138 25.6005
R4974 VDD.n140 VDD.n139 25.6005
R4975 VDD.n142 VDD.n140 25.6005
R4976 VDD.n143 VDD.n142 25.6005
R4977 VDD.n144 VDD.n143 25.6005
R4978 VDD.n145 VDD.n144 25.6005
R4979 VDD.n147 VDD.n145 25.6005
R4980 VDD.n148 VDD.n147 25.6005
R4981 VDD.n149 VDD.n148 25.6005
R4982 VDD.n150 VDD.n149 25.6005
R4983 VDD.n152 VDD.n150 25.6005
R4984 VDD.n153 VDD.n152 25.6005
R4985 VDD.n154 VDD.n153 25.6005
R4986 VDD.n155 VDD.n154 25.6005
R4987 VDD.n157 VDD.n155 25.6005
R4988 VDD.n158 VDD.n157 25.6005
R4989 VDD.n159 VDD.n158 25.6005
R4990 VDD.n160 VDD.n159 25.6005
R4991 VDD.n162 VDD.n160 25.6005
R4992 VDD.n163 VDD.n162 25.6005
R4993 VDD.n164 VDD.n163 25.6005
R4994 VDD.n83 VDD.n72 25.6005
R4995 VDD.n73 VDD.n72 25.6005
R4996 VDD.n76 VDD.n73 25.6005
R4997 VDD.n76 VDD.n48 25.6005
R4998 VDD.n303 VDD.n48 25.6005
R4999 VDD.n303 VDD.n302 25.6005
R5000 VDD.n52 VDD.n50 25.6005
R5001 VDD.n295 VDD.n52 25.6005
R5002 VDD.n295 VDD.n294 25.6005
R5003 VDD.n294 VDD.n293 25.6005
R5004 VDD.n293 VDD.n54 25.6005
R5005 VDD.n288 VDD.n287 25.6005
R5006 VDD.n287 VDD.n286 25.6005
R5007 VDD.n286 VDD.n57 25.6005
R5008 VDD.n281 VDD.n57 25.6005
R5009 VDD.n281 VDD.n280 25.6005
R5010 VDD.n280 VDD.n279 25.6005
R5011 VDD.n274 VDD.n60 25.6005
R5012 VDD.n274 VDD.n273 25.6005
R5013 VDD.n273 VDD.n272 25.6005
R5014 VDD.n272 VDD.n63 25.6005
R5015 VDD.n267 VDD.n63 25.6005
R5016 VDD.n349 VDD.t30 14.2851
R5017 VDD.n304 VDD.n303 11.5194
R5018 VDD.n263 VDD.t29 4.98619
R5019 VDD.n217 VDD.t43 4.98619
R5020 VDD.n257 VDD.t34 4.0797
R5021 VDD.n223 VDD.t2 4.0797
R5022 VDD.n323 VDD.n321 3.35217
R5023 VDD.n29 VDD.n27 3.35217
R5024 VDD.t3 VDD.n255 3.17321
R5025 VDD.n225 VDD.t7 3.17321
R5026 VDD.n4 VDD.n2 3.06997
R5027 VDD VDD.n354 2.80499
R5028 VDD.n341 VDD.n340 2.73818
R5029 VDD.n47 VDD.n46 2.73818
R5030 VDD.n351 VDD.n350 2.45598
R5031 VDD.n249 VDD.t22 2.26672
R5032 VDD.n231 VDD.t5 2.26672
R5033 VDD.n352 VDD.n341 2.07758
R5034 VDD.n354 VDD.n10 1.76955
R5035 VDD.n352 VDD.n351 1.63948
R5036 VDD.n304 VDD.n47 1.485
R5037 VDD.t17 VDD.n247 1.36023
R5038 VDD.n233 VDD.t11 1.36023
R5039 VDD.n353 VDD.n352 0.9725
R5040 VDD.n10 VDD.n8 0.61449
R5041 VDD.n8 VDD.n6 0.61449
R5042 VDD.n6 VDD.n4 0.61449
R5043 VDD.n351 VDD.n348 0.61449
R5044 VDD.n348 VDD.n346 0.61449
R5045 VDD.n346 VDD.n344 0.61449
R5046 VDD.n341 VDD.n323 0.61449
R5047 VDD.n47 VDD.n29 0.61449
R5048 VDD.n353 VDD.n304 0.590956
R5049 VDD.n354 VDD.n353 0.4865
R5050 VDD.n241 VDD.t0 0.453744
R5051 VDD.n239 VDD.t14 0.453744
R5052 VDD.n316 VDD.n307 0.38373
R5053 VDD.n311 VDD.n306 0.38373
R5054 VDD.n330 VDD.n329 0.38373
R5055 VDD.n336 VDD.n325 0.38373
R5056 VDD.n22 VDD.n21 0.383729
R5057 VDD.n15 VDD.n12 0.383729
R5058 VDD.n35 VDD.n33 0.383729
R5059 VDD.n42 VDD.n41 0.383729
R5060 VDD.n315 VDD.n308 0.338735
R5061 VDD.n308 VDD.n305 0.338735
R5062 VDD.n321 VDD.n305 0.338735
R5063 VDD.n335 VDD.n326 0.338735
R5064 VDD.n335 VDD.n324 0.338735
R5065 VDD.n340 VDD.n324 0.338735
R5066 VDD.n17 VDD.n13 0.338735
R5067 VDD.n17 VDD.n11 0.338735
R5068 VDD.n27 VDD.n11 0.338735
R5069 VDD.n36 VDD.n31 0.338735
R5070 VDD.n31 VDD.n30 0.338735
R5071 VDD.n46 VDD.n30 0.338735
R5072 VDD.n315 VDD.n314 0.285826
R5073 VDD.n309 VDD.n308 0.285826
R5074 VDD.n327 VDD.n326 0.285826
R5075 VDD.n335 VDD.n334 0.285826
R5076 VDD.n20 VDD.n13 0.285826
R5077 VDD.n18 VDD.n17 0.285826
R5078 VDD.n37 VDD.n36 0.285826
R5079 VDD.n39 VDD.n31 0.285826
R5080 VDD.n311 VDD.n310 0.188
R5081 VDD.n312 VDD.n311 0.188
R5082 VDD.n312 VDD.n307 0.188
R5083 VDD.n313 VDD.n309 0.188
R5084 VDD.n314 VDD.n313 0.188
R5085 VDD.n331 VDD.n330 0.188
R5086 VDD.n331 VDD.n325 0.188
R5087 VDD.n333 VDD.n325 0.188
R5088 VDD.n332 VDD.n327 0.188
R5089 VDD.n334 VDD.n332 0.188
R5090 VDD.n19 VDD.n18 0.188
R5091 VDD.n20 VDD.n19 0.188
R5092 VDD.n16 VDD.n15 0.188
R5093 VDD.n15 VDD.n14 0.188
R5094 VDD.n21 VDD.n14 0.188
R5095 VDD.n38 VDD.n37 0.188
R5096 VDD.n39 VDD.n38 0.188
R5097 VDD.n33 VDD.n32 0.188
R5098 VDD.n41 VDD.n32 0.188
R5099 VDD.n41 VDD.n40 0.188
R5100 VDD.n22 VDD.n13 0.0984044
R5101 VDD.n17 VDD.n12 0.0984044
R5102 VDD.n36 VDD.n35 0.0984044
R5103 VDD.n42 VDD.n31 0.0984044
R5104 VDD.n308 VDD.n306 0.0984028
R5105 VDD.n316 VDD.n315 0.0984028
R5106 VDD.n336 VDD.n335 0.0984028
R5107 VDD.n329 VDD.n326 0.0984028
R5108 VDD.n2 VDD.n1 0.0802101
R5109 a_6092_17969.n83 a_6092_17969.t25 260.486
R5110 a_6092_17969.n66 a_6092_17969.t27 260.486
R5111 a_6092_17969.n83 a_6092_17969.t21 260.111
R5112 a_6092_17969.n84 a_6092_17969.t32 260.111
R5113 a_6092_17969.n82 a_6092_17969.t23 260.111
R5114 a_6092_17969.n81 a_6092_17969.t24 260.111
R5115 a_6092_17969.n80 a_6092_17969.t34 260.111
R5116 a_6092_17969.n79 a_6092_17969.t31 260.111
R5117 a_6092_17969.n78 a_6092_17969.t22 260.111
R5118 a_6092_17969.n77 a_6092_17969.t33 260.111
R5119 a_6092_17969.n74 a_6092_17969.t19 260.111
R5120 a_6092_17969.n73 a_6092_17969.t30 260.111
R5121 a_6092_17969.n72 a_6092_17969.t26 260.111
R5122 a_6092_17969.n71 a_6092_17969.t18 260.111
R5123 a_6092_17969.n70 a_6092_17969.t28 260.111
R5124 a_6092_17969.n69 a_6092_17969.t29 260.111
R5125 a_6092_17969.n67 a_6092_17969.t20 260.111
R5126 a_6092_17969.n66 a_6092_17969.t35 260.111
R5127 a_6092_17969.n86 a_6092_17969.n85 203.843
R5128 a_6092_17969.n68 a_6092_17969.n65 203.843
R5129 a_6092_17969.n57 a_6092_17969.n39 185
R5130 a_6092_17969.n57 a_6092_17969.n38 185
R5131 a_6092_17969.n57 a_6092_17969.n37 185
R5132 a_6092_17969.n57 a_6092_17969.n36 185
R5133 a_6092_17969.n57 a_6092_17969.n35 185
R5134 a_6092_17969.n57 a_6092_17969.n34 185
R5135 a_6092_17969.n57 a_6092_17969.n33 185
R5136 a_6092_17969.n26 a_6092_17969.n8 185
R5137 a_6092_17969.n26 a_6092_17969.n7 185
R5138 a_6092_17969.n26 a_6092_17969.n6 185
R5139 a_6092_17969.n26 a_6092_17969.n5 185
R5140 a_6092_17969.n26 a_6092_17969.n4 185
R5141 a_6092_17969.n26 a_6092_17969.n3 185
R5142 a_6092_17969.n26 a_6092_17969.n2 185
R5143 a_6092_17969.n41 a_6092_17969.t7 130.75
R5144 a_6092_17969.n10 a_6092_17969.t5 130.75
R5145 a_6092_17969.n41 a_6092_17969.t9 91.3557
R5146 a_6092_17969.n10 a_6092_17969.t6 91.3557
R5147 a_6092_17969.n58 a_6092_17969.n57 86.5152
R5148 a_6092_17969.n27 a_6092_17969.n26 86.5152
R5149 a_6092_17969.n56 a_6092_17969.n40 30.3012
R5150 a_6092_17969.n25 a_6092_17969.n9 30.3012
R5151 a_6092_17969.n65 a_6092_17969.t2 28.5655
R5152 a_6092_17969.n65 a_6092_17969.t1 28.5655
R5153 a_6092_17969.t3 a_6092_17969.n86 28.5655
R5154 a_6092_17969.n86 a_6092_17969.t0 28.5655
R5155 a_6092_17969.n33 a_6092_17969.n32 24.8476
R5156 a_6092_17969.n2 a_6092_17969.n1 24.8476
R5157 a_6092_17969.n42 a_6092_17969.n34 23.3417
R5158 a_6092_17969.n11 a_6092_17969.n3 23.3417
R5159 a_6092_17969.n59 a_6092_17969.n58 22.0256
R5160 a_6092_17969.n28 a_6092_17969.n27 22.0256
R5161 a_6092_17969.n44 a_6092_17969.n35 21.8358
R5162 a_6092_17969.n13 a_6092_17969.n4 21.8358
R5163 a_6092_17969.n46 a_6092_17969.n36 20.3299
R5164 a_6092_17969.n15 a_6092_17969.n5 20.3299
R5165 a_6092_17969.n48 a_6092_17969.n37 18.824
R5166 a_6092_17969.n17 a_6092_17969.n6 18.824
R5167 a_6092_17969.n50 a_6092_17969.n38 17.3181
R5168 a_6092_17969.n19 a_6092_17969.n7 17.3181
R5169 a_6092_17969.n57 a_6092_17969.n56 16.3559
R5170 a_6092_17969.n26 a_6092_17969.n25 16.3559
R5171 a_6092_17969.n52 a_6092_17969.n39 15.8123
R5172 a_6092_17969.n21 a_6092_17969.n8 15.8123
R5173 a_6092_17969.n62 a_6092_17969.n61 14.6052
R5174 a_6092_17969.n64 a_6092_17969.n63 14.6052
R5175 a_6092_17969.n30 a_6092_17969.n29 14.377
R5176 a_6092_17969.n58 a_6092_17969.n32 12.7256
R5177 a_6092_17969.n27 a_6092_17969.n1 12.7256
R5178 a_6092_17969.n62 a_6092_17969.n60 11.5586
R5179 a_6092_17969.n40 a_6092_17969.n39 11.2946
R5180 a_6092_17969.n9 a_6092_17969.n8 11.2946
R5181 a_6092_17969.n75 a_6092_17969.t11 10.742
R5182 a_6092_17969.n52 a_6092_17969.n38 9.78874
R5183 a_6092_17969.n21 a_6092_17969.n7 9.78874
R5184 a_6092_17969.n32 a_6092_17969.n31 9.3005
R5185 a_6092_17969.n43 a_6092_17969.n42 9.3005
R5186 a_6092_17969.n45 a_6092_17969.n44 9.3005
R5187 a_6092_17969.n47 a_6092_17969.n46 9.3005
R5188 a_6092_17969.n49 a_6092_17969.n48 9.3005
R5189 a_6092_17969.n51 a_6092_17969.n50 9.3005
R5190 a_6092_17969.n53 a_6092_17969.n52 9.3005
R5191 a_6092_17969.n54 a_6092_17969.n40 9.3005
R5192 a_6092_17969.n1 a_6092_17969.n0 9.3005
R5193 a_6092_17969.n12 a_6092_17969.n11 9.3005
R5194 a_6092_17969.n14 a_6092_17969.n13 9.3005
R5195 a_6092_17969.n16 a_6092_17969.n15 9.3005
R5196 a_6092_17969.n18 a_6092_17969.n17 9.3005
R5197 a_6092_17969.n20 a_6092_17969.n19 9.3005
R5198 a_6092_17969.n22 a_6092_17969.n21 9.3005
R5199 a_6092_17969.n23 a_6092_17969.n9 9.3005
R5200 a_6092_17969.n76 a_6092_17969.n64 8.9511
R5201 a_6092_17969.n50 a_6092_17969.n37 8.28285
R5202 a_6092_17969.n19 a_6092_17969.n6 8.28285
R5203 a_6092_17969.n48 a_6092_17969.n36 6.77697
R5204 a_6092_17969.n17 a_6092_17969.n5 6.77697
R5205 a_6092_17969.n30 a_6092_17969.n28 6.19091
R5206 a_6092_17969.n46 a_6092_17969.n35 5.27109
R5207 a_6092_17969.n15 a_6092_17969.n4 5.27109
R5208 a_6092_17969.n44 a_6092_17969.n34 3.76521
R5209 a_6092_17969.n13 a_6092_17969.n3 3.76521
R5210 a_6092_17969.n60 a_6092_17969.n59 3.31388
R5211 a_6092_17969.n64 a_6092_17969.n62 2.87753
R5212 a_6092_17969.n75 a_6092_17969.n74 2.58895
R5213 a_6092_17969.n61 a_6092_17969.t12 2.48621
R5214 a_6092_17969.n61 a_6092_17969.t4 2.48621
R5215 a_6092_17969.n63 a_6092_17969.t17 2.48621
R5216 a_6092_17969.n63 a_6092_17969.t14 2.48621
R5217 a_6092_17969.n57 a_6092_17969.t15 2.48621
R5218 a_6092_17969.n57 a_6092_17969.t8 2.48621
R5219 a_6092_17969.n26 a_6092_17969.t6 2.48621
R5220 a_6092_17969.n26 a_6092_17969.t16 2.48621
R5221 a_6092_17969.n29 a_6092_17969.t13 2.48621
R5222 a_6092_17969.n29 a_6092_17969.t10 2.48621
R5223 a_6092_17969.n56 a_6092_17969.n55 2.36936
R5224 a_6092_17969.n25 a_6092_17969.n24 2.36936
R5225 a_6092_17969.n60 a_6092_17969.n30 2.30287
R5226 a_6092_17969.n42 a_6092_17969.n33 2.25932
R5227 a_6092_17969.n11 a_6092_17969.n2 2.25932
R5228 a_6092_17969.n76 a_6092_17969.n75 2.09432
R5229 a_6092_17969.n77 a_6092_17969.n76 1.78612
R5230 a_6092_17969.n67 a_6092_17969.n66 0.3755
R5231 a_6092_17969.n70 a_6092_17969.n69 0.3755
R5232 a_6092_17969.n71 a_6092_17969.n70 0.3755
R5233 a_6092_17969.n72 a_6092_17969.n71 0.3755
R5234 a_6092_17969.n73 a_6092_17969.n72 0.3755
R5235 a_6092_17969.n74 a_6092_17969.n73 0.3755
R5236 a_6092_17969.n78 a_6092_17969.n77 0.3755
R5237 a_6092_17969.n79 a_6092_17969.n78 0.3755
R5238 a_6092_17969.n80 a_6092_17969.n79 0.3755
R5239 a_6092_17969.n81 a_6092_17969.n80 0.3755
R5240 a_6092_17969.n82 a_6092_17969.n81 0.3755
R5241 a_6092_17969.n84 a_6092_17969.n83 0.3755
R5242 a_6092_17969.n55 a_6092_17969.n41 0.320353
R5243 a_6092_17969.n24 a_6092_17969.n10 0.320353
R5244 a_6092_17969.n55 a_6092_17969.n54 0.196152
R5245 a_6092_17969.n54 a_6092_17969.n53 0.196152
R5246 a_6092_17969.n53 a_6092_17969.n51 0.196152
R5247 a_6092_17969.n51 a_6092_17969.n49 0.196152
R5248 a_6092_17969.n49 a_6092_17969.n47 0.196152
R5249 a_6092_17969.n47 a_6092_17969.n45 0.196152
R5250 a_6092_17969.n45 a_6092_17969.n43 0.196152
R5251 a_6092_17969.n43 a_6092_17969.n31 0.196152
R5252 a_6092_17969.n59 a_6092_17969.n31 0.196152
R5253 a_6092_17969.n24 a_6092_17969.n23 0.196152
R5254 a_6092_17969.n23 a_6092_17969.n22 0.196152
R5255 a_6092_17969.n22 a_6092_17969.n20 0.196152
R5256 a_6092_17969.n20 a_6092_17969.n18 0.196152
R5257 a_6092_17969.n18 a_6092_17969.n16 0.196152
R5258 a_6092_17969.n16 a_6092_17969.n14 0.196152
R5259 a_6092_17969.n14 a_6092_17969.n12 0.196152
R5260 a_6092_17969.n12 a_6092_17969.n0 0.196152
R5261 a_6092_17969.n28 a_6092_17969.n0 0.196152
R5262 a_6092_17969.n68 a_6092_17969.n67 0.188
R5263 a_6092_17969.n69 a_6092_17969.n68 0.188
R5264 a_6092_17969.n85 a_6092_17969.n82 0.188
R5265 a_6092_17969.n85 a_6092_17969.n84 0.188
R5266 VOUT.n52 VOUT.t6 260.298
R5267 VOUT.t0 VOUT.n52 260.298
R5268 VOUT.t6 VOUT.n47 260.298
R5269 VOUT.t9 VOUT.n13 260.298
R5270 VOUT.n13 VOUT.t4 260.298
R5271 VOUT.t4 VOUT.n8 260.298
R5272 VOUT.n53 VOUT.t0 260.111
R5273 VOUT.n14 VOUT.t9 260.111
R5274 VOUT.n51 VOUT.t8 232.03
R5275 VOUT.n12 VOUT.t5 232.03
R5276 VOUT.n2 VOUT.n0 206.708
R5277 VOUT.n56 VOUT.n55 206.094
R5278 VOUT.n58 VOUT.n57 206.094
R5279 VOUT.n60 VOUT.n59 206.094
R5280 VOUT.n62 VOUT.n61 206.094
R5281 VOUT.n2 VOUT.n1 206.094
R5282 VOUT.n4 VOUT.n3 206.094
R5283 VOUT.n6 VOUT.n5 206.094
R5284 VOUT.n48 VOUT.n46 203.03
R5285 VOUT.n50 VOUT.n49 203.03
R5286 VOUT.n11 VOUT.n10 203.03
R5287 VOUT.n9 VOUT.n7 203.03
R5288 VOUT.n43 VOUT.n42 185
R5289 VOUT.n43 VOUT.n25 185
R5290 VOUT.n43 VOUT.n24 185
R5291 VOUT.n43 VOUT.n23 185
R5292 VOUT.n43 VOUT.n22 185
R5293 VOUT.n43 VOUT.n21 185
R5294 VOUT.n43 VOUT.n20 185
R5295 VOUT.n26 VOUT.t2 130.75
R5296 VOUT.n26 VOUT.t3 91.3557
R5297 VOUT.n44 VOUT.n43 86.5152
R5298 VOUT.n28 VOUT.n19 30.3012
R5299 VOUT.n63 VOUT.n45 29.1537
R5300 VOUT.n48 VOUT.t21 28.5655
R5301 VOUT.t1 VOUT.n48 28.5655
R5302 VOUT.n49 VOUT.t1 28.5655
R5303 VOUT.n49 VOUT.t7 28.5655
R5304 VOUT.n55 VOUT.t14 28.5655
R5305 VOUT.n55 VOUT.t25 28.5655
R5306 VOUT.n57 VOUT.t22 28.5655
R5307 VOUT.n57 VOUT.t23 28.5655
R5308 VOUT.n59 VOUT.t15 28.5655
R5309 VOUT.n59 VOUT.t12 28.5655
R5310 VOUT.n61 VOUT.t13 28.5655
R5311 VOUT.n61 VOUT.t24 28.5655
R5312 VOUT.n0 VOUT.t16 28.5655
R5313 VOUT.n0 VOUT.t27 28.5655
R5314 VOUT.n1 VOUT.t28 28.5655
R5315 VOUT.n1 VOUT.t20 28.5655
R5316 VOUT.n3 VOUT.t17 28.5655
R5317 VOUT.n3 VOUT.t18 28.5655
R5318 VOUT.n5 VOUT.t11 28.5655
R5319 VOUT.n5 VOUT.t26 28.5655
R5320 VOUT.n10 VOUT.t5 28.5655
R5321 VOUT.n10 VOUT.t10 28.5655
R5322 VOUT.t10 VOUT.n9 28.5655
R5323 VOUT.n9 VOUT.t19 28.5655
R5324 VOUT.n42 VOUT.n18 24.8476
R5325 VOUT.n41 VOUT.n25 23.3417
R5326 VOUT.n45 VOUT.n44 22.0256
R5327 VOUT.n38 VOUT.n24 21.8358
R5328 VOUT.n36 VOUT.n23 20.3299
R5329 VOUT.n34 VOUT.n22 18.824
R5330 VOUT.n32 VOUT.n21 17.3181
R5331 VOUT.n43 VOUT.n19 16.3559
R5332 VOUT.n30 VOUT.n20 15.8123
R5333 VOUT.n44 VOUT.n18 12.7256
R5334 VOUT.n28 VOUT.n20 11.2946
R5335 VOUT.n30 VOUT.n21 9.78874
R5336 VOUT.n18 VOUT.n17 9.3005
R5337 VOUT.n41 VOUT.n40 9.3005
R5338 VOUT.n39 VOUT.n38 9.3005
R5339 VOUT.n37 VOUT.n36 9.3005
R5340 VOUT.n35 VOUT.n34 9.3005
R5341 VOUT.n33 VOUT.n32 9.3005
R5342 VOUT.n31 VOUT.n30 9.3005
R5343 VOUT.n29 VOUT.n28 9.3005
R5344 VOUT.n32 VOUT.n22 8.28285
R5345 VOUT.n65 VOUT.n64 8.02834
R5346 VOUT.n34 VOUT.n23 6.77697
R5347 VOUT.n36 VOUT.n24 5.27109
R5348 VOUT.n38 VOUT.n25 3.76521
R5349 VOUT.n63 VOUT.n62 3.22728
R5350 VOUT.n56 VOUT.n54 3.17011
R5351 VOUT.n16 VOUT.n15 2.55612
R5352 VOUT.n43 VOUT.t3 2.48621
R5353 VOUT.n43 VOUT.t30 2.48621
R5354 VOUT.n27 VOUT.n19 2.36936
R5355 VOUT.n42 VOUT.n41 2.25932
R5356 VOUT.n64 VOUT.n16 2.22267
R5357 VOUT.n64 VOUT 0.774914
R5358 VOUT.n62 VOUT.n60 0.61449
R5359 VOUT.n60 VOUT.n58 0.61449
R5360 VOUT.n58 VOUT.n56 0.61449
R5361 VOUT.n16 VOUT.n6 0.61449
R5362 VOUT.n6 VOUT.n4 0.61449
R5363 VOUT.n4 VOUT.n2 0.61449
R5364 VOUT.n51 VOUT.n46 0.43664
R5365 VOUT.n12 VOUT.n7 0.436638
R5366 VOUT.n15 VOUT.n7 0.38373
R5367 VOUT.n11 VOUT.n8 0.38373
R5368 VOUT.n54 VOUT.n46 0.383729
R5369 VOUT.n50 VOUT.n47 0.383729
R5370 VOUT.n27 VOUT.n26 0.320353
R5371 VOUT.n52 VOUT.n51 0.285826
R5372 VOUT.n13 VOUT.n12 0.285826
R5373 VOUT.n45 VOUT.n17 0.196152
R5374 VOUT.n40 VOUT.n17 0.196152
R5375 VOUT.n40 VOUT.n39 0.196152
R5376 VOUT.n39 VOUT.n37 0.196152
R5377 VOUT.n37 VOUT.n35 0.196152
R5378 VOUT.n35 VOUT.n33 0.196152
R5379 VOUT.n33 VOUT.n31 0.196152
R5380 VOUT.n31 VOUT.n29 0.196152
R5381 VOUT.n29 VOUT.n27 0.196152
R5382 VOUT.n54 VOUT.n53 0.188
R5383 VOUT.n53 VOUT.n47 0.188
R5384 VOUT.n14 VOUT.n8 0.188
R5385 VOUT.n15 VOUT.n14 0.188
R5386 VOUT VOUT.n65 0.185987
R5387 VOUT VOUT.n63 0.113781
R5388 VOUT.n51 VOUT.n50 0.0984044
R5389 VOUT.n12 VOUT.n11 0.0984028
R5390 VOUT.n65 VOUT.t29 0.0409532
R5391 VP.n0 VP.t7 263.647
R5392 VP.n3 VP.t5 262.863
R5393 VP.n2 VP.t6 262.498
R5394 VP.n0 VP.t2 261.709
R5395 VP.n1 VP.t4 261.709
R5396 VP.n3 VP.t1 261.584
R5397 VP.n4 VP.t3 261.584
R5398 VP.n5 VP.t0 261.433
R5399 VP.n6 VP.n2 8.91142
R5400 VP VP.n6 3.01373
R5401 VP.n1 VP.n0 1.72698
R5402 VP.n6 VP.n5 1.52193
R5403 VP.n5 VP.n4 1.4312
R5404 VP.n4 VP.n3 1.16675
R5405 VP.n2 VP.n1 1.14999
R5406 a_6105_7756.n23 a_6105_7756.n1 185
R5407 a_6105_7756.n25 a_6105_7756.n1 185
R5408 a_6105_7756.n4 a_6105_7756.n1 185
R5409 a_6105_7756.n30 a_6105_7756.n1 185
R5410 a_6105_7756.n32 a_6105_7756.n1 185
R5411 a_6105_7756.n2 a_6105_7756.n1 185
R5412 a_6105_7756.n37 a_6105_7756.n1 185
R5413 a_6105_7756.t2 a_6105_7756.n42 180.167
R5414 a_6105_7756.t2 a_6105_7756.n42 180.167
R5415 a_6105_7756.n41 a_6105_7756.t0 130.75
R5416 a_6105_7756.n6 a_6105_7756.n1 86.5152
R5417 a_6105_7756.n39 a_6105_7756.n38 30.3012
R5418 a_6105_7756.n23 a_6105_7756.n22 24.8476
R5419 a_6105_7756.n25 a_6105_7756.n24 23.3417
R5420 a_6105_7756.n20 a_6105_7756.n6 22.0256
R5421 a_6105_7756.n26 a_6105_7756.n4 21.8358
R5422 a_6105_7756.n30 a_6105_7756.n29 20.3299
R5423 a_6105_7756.n32 a_6105_7756.n31 18.824
R5424 a_6105_7756.n33 a_6105_7756.n2 17.3181
R5425 a_6105_7756.n39 a_6105_7756.n1 16.3559
R5426 a_6105_7756.n37 a_6105_7756.n36 15.8123
R5427 a_6105_7756.n22 a_6105_7756.n6 12.7256
R5428 a_6105_7756.n9 a_6105_7756.n7 11.493
R5429 a_6105_7756.n16 a_6105_7756.n14 11.493
R5430 a_6105_7756.n17 a_6105_7756.n12 11.493
R5431 a_6105_7756.n18 a_6105_7756.n10 11.493
R5432 a_6105_7756.n9 a_6105_7756.n8 11.4929
R5433 a_6105_7756.n16 a_6105_7756.n15 11.4929
R5434 a_6105_7756.n17 a_6105_7756.n13 11.4929
R5435 a_6105_7756.n18 a_6105_7756.n11 11.4929
R5436 a_6105_7756.n38 a_6105_7756.n37 11.2946
R5437 a_6105_7756.n19 a_6105_7756.n18 9.83015
R5438 a_6105_7756.n19 a_6105_7756.n9 9.83015
R5439 a_6105_7756.n36 a_6105_7756.n2 9.78874
R5440 a_6105_7756.n22 a_6105_7756.n21 9.3005
R5441 a_6105_7756.n24 a_6105_7756.n5 9.3005
R5442 a_6105_7756.n27 a_6105_7756.n26 9.3005
R5443 a_6105_7756.n29 a_6105_7756.n28 9.3005
R5444 a_6105_7756.n31 a_6105_7756.n3 9.3005
R5445 a_6105_7756.n34 a_6105_7756.n33 9.3005
R5446 a_6105_7756.n36 a_6105_7756.n35 9.3005
R5447 a_6105_7756.n38 a_6105_7756.n0 9.3005
R5448 a_6105_7756.n33 a_6105_7756.n32 8.28285
R5449 a_6105_7756.n31 a_6105_7756.n30 6.77697
R5450 a_6105_7756.n20 a_6105_7756.n19 6.3915
R5451 a_6105_7756.n29 a_6105_7756.n4 5.27109
R5452 a_6105_7756.n26 a_6105_7756.n25 3.76521
R5453 a_6105_7756.n1 a_6105_7756.t8 2.48621
R5454 a_6105_7756.n1 a_6105_7756.t1 2.48621
R5455 a_6105_7756.n8 a_6105_7756.t16 2.48621
R5456 a_6105_7756.n8 a_6105_7756.t17 2.48621
R5457 a_6105_7756.n7 a_6105_7756.t19 2.48621
R5458 a_6105_7756.n7 a_6105_7756.t10 2.48621
R5459 a_6105_7756.n15 a_6105_7756.t6 2.48621
R5460 a_6105_7756.n15 a_6105_7756.t13 2.48621
R5461 a_6105_7756.n14 a_6105_7756.t12 2.48621
R5462 a_6105_7756.n14 a_6105_7756.t7 2.48621
R5463 a_6105_7756.n13 a_6105_7756.t15 2.48621
R5464 a_6105_7756.n13 a_6105_7756.t3 2.48621
R5465 a_6105_7756.n12 a_6105_7756.t4 2.48621
R5466 a_6105_7756.n12 a_6105_7756.t14 2.48621
R5467 a_6105_7756.n11 a_6105_7756.t5 2.48621
R5468 a_6105_7756.n11 a_6105_7756.t11 2.48621
R5469 a_6105_7756.n10 a_6105_7756.t9 2.48621
R5470 a_6105_7756.n10 a_6105_7756.t18 2.48621
R5471 a_6105_7756.n40 a_6105_7756.n39 2.36936
R5472 a_6105_7756.n24 a_6105_7756.n23 2.25932
R5473 a_6105_7756.n42 a_6105_7756.n41 1.27148
R5474 a_6105_7756.n16 a_6105_7756.n9 1.15229
R5475 a_6105_7756.n17 a_6105_7756.n16 1.15229
R5476 a_6105_7756.n18 a_6105_7756.n17 1.15229
R5477 a_6105_7756.n41 a_6105_7756.n40 0.320353
R5478 a_6105_7756.n21 a_6105_7756.n20 0.196152
R5479 a_6105_7756.n21 a_6105_7756.n5 0.196152
R5480 a_6105_7756.n27 a_6105_7756.n5 0.196152
R5481 a_6105_7756.n28 a_6105_7756.n27 0.196152
R5482 a_6105_7756.n28 a_6105_7756.n3 0.196152
R5483 a_6105_7756.n34 a_6105_7756.n3 0.196152
R5484 a_6105_7756.n35 a_6105_7756.n34 0.196152
R5485 a_6105_7756.n35 a_6105_7756.n0 0.196152
R5486 a_6105_7756.n40 a_6105_7756.n0 0.196152
R5487 a_6423_5719.n39 a_6423_5719.n4 185
R5488 a_6423_5719.n39 a_6423_5719.n6 185
R5489 a_6423_5719.n39 a_6423_5719.n3 185
R5490 a_6423_5719.n39 a_6423_5719.n7 185
R5491 a_6423_5719.n39 a_6423_5719.n2 185
R5492 a_6423_5719.n39 a_6423_5719.n8 185
R5493 a_6423_5719.n39 a_6423_5719.n1 185
R5494 a_6423_5719.n0 a_6423_5719.t0 130.75
R5495 a_6423_5719.t1 a_6423_5719.n0 91.3557
R5496 a_6423_5719.n39 a_6423_5719.n5 86.5152
R5497 a_6423_5719.n38 a_6423_5719.n37 30.3012
R5498 a_6423_5719.n12 a_6423_5719.n10 29.1073
R5499 a_6423_5719.n12 a_6423_5719.n11 27.9576
R5500 a_6423_5719.n14 a_6423_5719.n13 27.9576
R5501 a_6423_5719.n16 a_6423_5719.n15 27.9576
R5502 a_6423_5719.n18 a_6423_5719.n17 27.9576
R5503 a_6423_5719.n20 a_6423_5719.n19 27.9576
R5504 a_6423_5719.n22 a_6423_5719.n4 24.8476
R5505 a_6423_5719.n24 a_6423_5719.n6 23.3417
R5506 a_6423_5719.n21 a_6423_5719.n5 22.0256
R5507 a_6423_5719.n26 a_6423_5719.n3 21.8358
R5508 a_6423_5719.n28 a_6423_5719.n7 20.3299
R5509 a_6423_5719.n30 a_6423_5719.n2 18.824
R5510 a_6423_5719.n32 a_6423_5719.n8 17.3181
R5511 a_6423_5719.n39 a_6423_5719.n38 16.3559
R5512 a_6423_5719.n34 a_6423_5719.n1 15.8123
R5513 a_6423_5719.n22 a_6423_5719.n5 12.7256
R5514 a_6423_5719.n37 a_6423_5719.n1 11.2946
R5515 a_6423_5719.n21 a_6423_5719.n20 10.9789
R5516 a_6423_5719.n34 a_6423_5719.n8 9.78874
R5517 a_6423_5719.n23 a_6423_5719.n22 9.3005
R5518 a_6423_5719.n25 a_6423_5719.n24 9.3005
R5519 a_6423_5719.n27 a_6423_5719.n26 9.3005
R5520 a_6423_5719.n29 a_6423_5719.n28 9.3005
R5521 a_6423_5719.n31 a_6423_5719.n30 9.3005
R5522 a_6423_5719.n33 a_6423_5719.n32 9.3005
R5523 a_6423_5719.n35 a_6423_5719.n34 9.3005
R5524 a_6423_5719.n37 a_6423_5719.n36 9.3005
R5525 a_6423_5719.n32 a_6423_5719.n2 8.28285
R5526 a_6423_5719.n30 a_6423_5719.n7 6.77697
R5527 a_6423_5719.n10 a_6423_5719.t7 5.8005
R5528 a_6423_5719.n10 a_6423_5719.t9 5.8005
R5529 a_6423_5719.n11 a_6423_5719.t8 5.8005
R5530 a_6423_5719.n11 a_6423_5719.t13 5.8005
R5531 a_6423_5719.n13 a_6423_5719.t4 5.8005
R5532 a_6423_5719.n13 a_6423_5719.t3 5.8005
R5533 a_6423_5719.n15 a_6423_5719.t11 5.8005
R5534 a_6423_5719.n15 a_6423_5719.t10 5.8005
R5535 a_6423_5719.n17 a_6423_5719.t2 5.8005
R5536 a_6423_5719.n17 a_6423_5719.t12 5.8005
R5537 a_6423_5719.n19 a_6423_5719.t5 5.8005
R5538 a_6423_5719.n19 a_6423_5719.t6 5.8005
R5539 a_6423_5719.n28 a_6423_5719.n3 5.27109
R5540 a_6423_5719.n26 a_6423_5719.n6 3.76521
R5541 a_6423_5719.t1 a_6423_5719.n39 2.48621
R5542 a_6423_5719.n39 a_6423_5719.t14 2.48621
R5543 a_6423_5719.n38 a_6423_5719.n9 2.36936
R5544 a_6423_5719.n16 a_6423_5719.n14 2.30199
R5545 a_6423_5719.n24 a_6423_5719.n4 2.25932
R5546 a_6423_5719.n20 a_6423_5719.n18 1.1502
R5547 a_6423_5719.n18 a_6423_5719.n16 1.1502
R5548 a_6423_5719.n14 a_6423_5719.n12 1.1502
R5549 a_6423_5719.n9 a_6423_5719.n0 0.320353
R5550 a_6423_5719.n23 a_6423_5719.n21 0.196152
R5551 a_6423_5719.n25 a_6423_5719.n23 0.196152
R5552 a_6423_5719.n27 a_6423_5719.n25 0.196152
R5553 a_6423_5719.n29 a_6423_5719.n27 0.196152
R5554 a_6423_5719.n31 a_6423_5719.n29 0.196152
R5555 a_6423_5719.n33 a_6423_5719.n31 0.196152
R5556 a_6423_5719.n35 a_6423_5719.n33 0.196152
R5557 a_6423_5719.n36 a_6423_5719.n35 0.196152
R5558 a_6423_5719.n36 a_6423_5719.n9 0.196152
R5559 VN.n0 VN.t6 263.647
R5560 VN.n3 VN.t1 262.863
R5561 VN.n2 VN.t7 262.498
R5562 VN.n1 VN.t0 261.709
R5563 VN.n0 VN.t3 261.709
R5564 VN.n4 VN.t2 261.584
R5565 VN.n3 VN.t4 261.584
R5566 VN.n5 VN.t5 261.433
R5567 VN.n6 VN.n2 8.91142
R5568 VN VN.n6 3.22767
R5569 VN.n1 VN.n0 1.72698
R5570 VN.n6 VN.n5 1.52193
R5571 VN.n5 VN.n4 1.4312
R5572 VN.n4 VN.n3 1.16675
R5573 VN.n2 VN.n1 1.14999
R5574 EN.n0 EN.t0 262.997
R5575 EN.n1 EN.t1 262.007
R5576 EN.n0 EN.t2 262.007
R5577 EN.n1 EN.n0 0.989232
R5578 EN EN.n1 0.359662
R5579 C1 C1.t0 16.6024
R5580 C1 C1.t1 0.00167066
R5581 IBIAS.n26 IBIAS.n25 185
R5582 IBIAS.n26 IBIAS.n8 185
R5583 IBIAS.n26 IBIAS.n7 185
R5584 IBIAS.n26 IBIAS.n6 185
R5585 IBIAS.n26 IBIAS.n5 185
R5586 IBIAS.n26 IBIAS.n4 185
R5587 IBIAS.n26 IBIAS.n3 185
R5588 IBIAS.n9 IBIAS.t1 130.75
R5589 IBIAS.n9 IBIAS.t2 91.3557
R5590 IBIAS.n27 IBIAS.n26 86.5152
R5591 IBIAS.n11 IBIAS.n2 30.3012
R5592 IBIAS.n25 IBIAS.n1 24.8476
R5593 IBIAS.n24 IBIAS.n8 23.3417
R5594 IBIAS.n28 IBIAS.n27 22.0256
R5595 IBIAS.n21 IBIAS.n7 21.8358
R5596 IBIAS.n19 IBIAS.n6 20.3299
R5597 IBIAS.n17 IBIAS.n5 18.824
R5598 IBIAS.n15 IBIAS.n4 17.3181
R5599 IBIAS.n26 IBIAS.n2 16.3559
R5600 IBIAS.n13 IBIAS.n3 15.8123
R5601 IBIAS.n27 IBIAS.n1 12.7256
R5602 IBIAS.n11 IBIAS.n3 11.2946
R5603 IBIAS.n13 IBIAS.n4 9.78874
R5604 IBIAS.n1 IBIAS.n0 9.3005
R5605 IBIAS.n24 IBIAS.n23 9.3005
R5606 IBIAS.n22 IBIAS.n21 9.3005
R5607 IBIAS.n20 IBIAS.n19 9.3005
R5608 IBIAS.n18 IBIAS.n17 9.3005
R5609 IBIAS.n16 IBIAS.n15 9.3005
R5610 IBIAS.n14 IBIAS.n13 9.3005
R5611 IBIAS.n12 IBIAS.n11 9.3005
R5612 IBIAS.n15 IBIAS.n5 8.28285
R5613 IBIAS IBIAS.n28 8.01267
R5614 IBIAS.n17 IBIAS.n6 6.77697
R5615 IBIAS.n19 IBIAS.n7 5.27109
R5616 IBIAS.n21 IBIAS.n8 3.76521
R5617 IBIAS.n26 IBIAS.t2 2.48621
R5618 IBIAS.n26 IBIAS.t0 2.48621
R5619 IBIAS.n10 IBIAS.n2 2.36936
R5620 IBIAS.n25 IBIAS.n24 2.25932
R5621 IBIAS.n10 IBIAS.n9 0.320353
R5622 IBIAS.n28 IBIAS.n0 0.196152
R5623 IBIAS.n23 IBIAS.n0 0.196152
R5624 IBIAS.n23 IBIAS.n22 0.196152
R5625 IBIAS.n22 IBIAS.n20 0.196152
R5626 IBIAS.n20 IBIAS.n18 0.196152
R5627 IBIAS.n18 IBIAS.n16 0.196152
R5628 IBIAS.n16 IBIAS.n14 0.196152
R5629 IBIAS.n14 IBIAS.n12 0.196152
R5630 IBIAS.n12 IBIAS.n10 0.196152
C6 IBIAS VSS 2.47026f
C7 EN VSS 2.86135f
C8 VP VSS 6.2001f
C9 VN VSS 6.16092f
C10 VOUT VSS 23.20691f
C11 VDD VSS 14.70285f
C12 C1 VSS 32.58249f $ **FLOATING
C13 C1.t0 VSS 0.23907f $ **FLOATING
C14 C1.t1 VSS 28.8988f $ **FLOATING
C15 VN.t6 VSS 1.34251f $ **FLOATING
C16 VN.t3 VSS 1.33868f $ **FLOATING
C17 VN.n0 VSS 1.18156f $ **FLOATING
C18 VN.t0 VSS 1.33868f $ **FLOATING
C19 VN.n1 VSS 0.59f $ **FLOATING
C20 VN.t7 VSS 1.33992f $ **FLOATING
C21 VN.n2 VSS 1.05074f $ **FLOATING
C22 VN.t2 VSS 1.33838f $ **FLOATING
C23 VN.t1 VSS 1.3415f $ **FLOATING
C24 VN.t4 VSS 1.33838f $ **FLOATING
C25 VN.n3 VSS 1.16738f $ **FLOATING
C26 VN.n4 VSS 0.55877f $ **FLOATING
C27 VN.t5 VSS 1.33817f $ **FLOATING
C28 VN.n5 VSS 0.57983f $ **FLOATING
C29 VN.n6 VSS 0.80581f $ **FLOATING
C30 a_6423_5719.t0 VSS 0.44262f $ **FLOATING
C31 a_6423_5719.n0 VSS 0.83924f $ **FLOATING
C32 a_6423_5719.t14 VSS 0.04451f $ **FLOATING
C33 a_6423_5719.n9 VSS 0.11938f $ **FLOATING
C34 a_6423_5719.t7 VSS 0.01907f $ **FLOATING
C35 a_6423_5719.t9 VSS 0.01907f $ **FLOATING
C36 a_6423_5719.n10 VSS 0.06586f $ **FLOATING
C37 a_6423_5719.t8 VSS 0.01907f $ **FLOATING
C38 a_6423_5719.t13 VSS 0.01907f $ **FLOATING
C39 a_6423_5719.n11 VSS 0.05604f $ **FLOATING
C40 a_6423_5719.n12 VSS 0.42796f $ **FLOATING
C41 a_6423_5719.t4 VSS 0.01907f $ **FLOATING
C42 a_6423_5719.t3 VSS 0.01907f $ **FLOATING
C43 a_6423_5719.n13 VSS 0.05604f $ **FLOATING
C44 a_6423_5719.n14 VSS 0.22079f $ **FLOATING
C45 a_6423_5719.t11 VSS 0.01907f $ **FLOATING
C46 a_6423_5719.t10 VSS 0.01907f $ **FLOATING
C47 a_6423_5719.n15 VSS 0.05604f $ **FLOATING
C48 a_6423_5719.n16 VSS 0.22079f $ **FLOATING
C49 a_6423_5719.t2 VSS 0.01907f $ **FLOATING
C50 a_6423_5719.t12 VSS 0.01907f $ **FLOATING
C51 a_6423_5719.n17 VSS 0.05604f $ **FLOATING
C52 a_6423_5719.n18 VSS 0.18912f $ **FLOATING
C53 a_6423_5719.t5 VSS 0.01907f $ **FLOATING
C54 a_6423_5719.t6 VSS 0.01907f $ **FLOATING
C55 a_6423_5719.n19 VSS 0.05604f $ **FLOATING
C56 a_6423_5719.n20 VSS 2.00961f $ **FLOATING
C57 a_6423_5719.n21 VSS 1.43678f $ **FLOATING
C58 a_6423_5719.n39 VSS 0.09522f $ **FLOATING
C59 a_6423_5719.t1 VSS 0.06801f $ **FLOATING
C60 a_6105_7756.n0 VSS 0.01462f $ **FLOATING
C61 a_6105_7756.t8 VSS 0.08962f $ **FLOATING
C62 a_6105_7756.t1 VSS 0.08962f $ **FLOATING
C63 a_6105_7756.n1 VSS 0.19173f $ **FLOATING
C64 a_6105_7756.n3 VSS 0.01462f $ **FLOATING
C65 a_6105_7756.n5 VSS 0.01462f $ **FLOATING
C66 a_6105_7756.t19 VSS 0.08962f $ **FLOATING
C67 a_6105_7756.t10 VSS 0.08962f $ **FLOATING
C68 a_6105_7756.n7 VSS 0.25639f $ **FLOATING
C69 a_6105_7756.t16 VSS 0.08962f $ **FLOATING
C70 a_6105_7756.t17 VSS 0.08962f $ **FLOATING
C71 a_6105_7756.n8 VSS 0.25641f $ **FLOATING
C72 a_6105_7756.n9 VSS 1.19281f $ **FLOATING
C73 a_6105_7756.t9 VSS 0.08962f $ **FLOATING
C74 a_6105_7756.t18 VSS 0.08962f $ **FLOATING
C75 a_6105_7756.n10 VSS 0.25639f $ **FLOATING
C76 a_6105_7756.t5 VSS 0.08962f $ **FLOATING
C77 a_6105_7756.t11 VSS 0.08962f $ **FLOATING
C78 a_6105_7756.n11 VSS 0.25641f $ **FLOATING
C79 a_6105_7756.t4 VSS 0.08962f $ **FLOATING
C80 a_6105_7756.t14 VSS 0.08962f $ **FLOATING
C81 a_6105_7756.n12 VSS 0.25639f $ **FLOATING
C82 a_6105_7756.t15 VSS 0.08962f $ **FLOATING
C83 a_6105_7756.t3 VSS 0.08962f $ **FLOATING
C84 a_6105_7756.n13 VSS 0.25641f $ **FLOATING
C85 a_6105_7756.t12 VSS 0.08962f $ **FLOATING
C86 a_6105_7756.t7 VSS 0.08962f $ **FLOATING
C87 a_6105_7756.n14 VSS 0.25639f $ **FLOATING
C88 a_6105_7756.t6 VSS 0.08962f $ **FLOATING
C89 a_6105_7756.t13 VSS 0.08962f $ **FLOATING
C90 a_6105_7756.n15 VSS 0.25641f $ **FLOATING
C91 a_6105_7756.n16 VSS 1.00758f $ **FLOATING
C92 a_6105_7756.n17 VSS 1.00758f $ **FLOATING
C93 a_6105_7756.n18 VSS 1.2082f $ **FLOATING
C94 a_6105_7756.n19 VSS 4.94247f $ **FLOATING
C95 a_6105_7756.n20 VSS 0.29278f $ **FLOATING
C96 a_6105_7756.n21 VSS 0.01462f $ **FLOATING
C97 a_6105_7756.n22 VSS 0.01005f $ **FLOATING
C98 a_6105_7756.n27 VSS 0.01462f $ **FLOATING
C99 a_6105_7756.n28 VSS 0.01462f $ **FLOATING
C100 a_6105_7756.n34 VSS 0.01462f $ **FLOATING
C101 a_6105_7756.n35 VSS 0.01462f $ **FLOATING
C102 a_6105_7756.n39 VSS 0.0121f $ **FLOATING
C103 a_6105_7756.n40 VSS 0.24038f $ **FLOATING
C104 a_6105_7756.t0 VSS 0.89127f $ **FLOATING
C105 a_6105_7756.n41 VSS 1.43629f $ **FLOATING
C106 a_6105_7756.n42 VSS 0.25721f $ **FLOATING
C107 a_6105_7756.t2 VSS 0.04375f $ **FLOATING
C108 VP.t7 VSS 1.33483f $ **FLOATING
C109 VP.t2 VSS 1.33103f $ **FLOATING
C110 VP.n0 VSS 1.17481f $ **FLOATING
C111 VP.t4 VSS 1.33103f $ **FLOATING
C112 VP.n1 VSS 0.58663f $ **FLOATING
C113 VP.t6 VSS 1.33226f $ **FLOATING
C114 VP.n2 VSS 1.04473f $ **FLOATING
C115 VP.t5 VSS 1.33383f $ **FLOATING
C116 VP.t1 VSS 1.33073f $ **FLOATING
C117 VP.n3 VSS 1.1607f $ **FLOATING
C118 VP.t3 VSS 1.33073f $ **FLOATING
C119 VP.n4 VSS 0.55557f $ **FLOATING
C120 VP.t0 VSS 1.33052f $ **FLOATING
C121 VP.n5 VSS 0.57652f $ **FLOATING
C122 VP.n6 VSS 0.7502f $ **FLOATING
C123 VOUT.t29 VSS 51.7429f $ **FLOATING
C124 VOUT.n0 VSS 0.01463f $ **FLOATING
C125 VOUT.n1 VSS 0.01418f $ **FLOATING
C126 VOUT.n2 VSS 0.25924f $ **FLOATING
C127 VOUT.n3 VSS 0.01418f $ **FLOATING
C128 VOUT.n4 VSS 0.10881f $ **FLOATING
C129 VOUT.n5 VSS 0.01418f $ **FLOATING
C130 VOUT.n6 VSS 0.10881f $ **FLOATING
C131 VOUT.n7 VSS 0.02994f $ **FLOATING
C132 VOUT.n8 VSS 0.03599f $ **FLOATING
C133 VOUT.t4 VSS 0.05403f $ **FLOATING
C134 VOUT.t5 VSS 0.02986f $ **FLOATING
C135 VOUT.n9 VSS 0.0132f $ **FLOATING
C136 VOUT.t10 VSS 0.01267f $ **FLOATING
C137 VOUT.n10 VSS 0.0132f $ **FLOATING
C138 VOUT.n11 VSS 0.01623f $ **FLOATING
C139 VOUT.n12 VSS 0.06468f $ **FLOATING
C140 VOUT.n13 VSS 0.05307f $ **FLOATING
C141 VOUT.t9 VSS 0.05401f $ **FLOATING
C142 VOUT.n14 VSS 0.02029f $ **FLOATING
C143 VOUT.n15 VSS 0.04325f $ **FLOATING
C144 VOUT.n16 VSS 0.08116f $ **FLOATING
C145 VOUT.t3 VSS 0.06775f $ **FLOATING
C146 VOUT.t2 VSS 0.44093f $ **FLOATING
C147 VOUT.n26 VSS 0.83605f $ **FLOATING
C148 VOUT.n27 VSS 0.11892f $ **FLOATING
C149 VOUT.t30 VSS 0.04434f $ **FLOATING
C150 VOUT.n43 VSS 0.09485f $ **FLOATING
C151 VOUT.n45 VSS 0.68892f $ **FLOATING
C152 VOUT.n46 VSS 0.02994f $ **FLOATING
C153 VOUT.n47 VSS 0.03599f $ **FLOATING
C154 VOUT.t6 VSS 0.05403f $ **FLOATING
C155 VOUT.t8 VSS 0.02353f $ **FLOATING
C156 VOUT.n48 VSS 0.0132f $ **FLOATING
C157 VOUT.t1 VSS 0.01267f $ **FLOATING
C158 VOUT.n49 VSS 0.0132f $ **FLOATING
C159 VOUT.n50 VSS 0.01623f $ **FLOATING
C160 VOUT.n51 VSS 0.06468f $ **FLOATING
C161 VOUT.n52 VSS 0.05307f $ **FLOATING
C162 VOUT.t0 VSS 0.05401f $ **FLOATING
C163 VOUT.n53 VSS 0.02029f $ **FLOATING
C164 VOUT.n54 VSS 0.05859f $ **FLOATING
C165 VOUT.n55 VSS 0.01418f $ **FLOATING
C166 VOUT.n56 VSS 0.17274f $ **FLOATING
C167 VOUT.n57 VSS 0.01418f $ **FLOATING
C168 VOUT.n58 VSS 0.10881f $ **FLOATING
C169 VOUT.n59 VSS 0.01418f $ **FLOATING
C170 VOUT.n60 VSS 0.10881f $ **FLOATING
C171 VOUT.n61 VSS 0.01418f $ **FLOATING
C172 VOUT.n62 VSS 0.23034f $ **FLOATING
C173 VOUT.n63 VSS 1.1168f $ **FLOATING
C174 VOUT.n64 VSS 0.83445f $ **FLOATING
C175 VOUT.n65 VSS 11.984f $ **FLOATING
C176 a_6092_17969.n0 VSS 0.0169f $ **FLOATING
C177 a_6092_17969.n1 VSS 0.01161f $ **FLOATING
C178 a_6092_17969.t6 VSS 0.15828f $ **FLOATING
C179 a_6092_17969.n9 VSS 0.01126f $ **FLOATING
C180 a_6092_17969.t5 VSS 1.03028f $ **FLOATING
C181 a_6092_17969.n10 VSS 1.97223f $ **FLOATING
C182 a_6092_17969.n12 VSS 0.0169f $ **FLOATING
C183 a_6092_17969.n14 VSS 0.0169f $ **FLOATING
C184 a_6092_17969.n16 VSS 0.0169f $ **FLOATING
C185 a_6092_17969.n18 VSS 0.0169f $ **FLOATING
C186 a_6092_17969.n20 VSS 0.0169f $ **FLOATING
C187 a_6092_17969.n22 VSS 0.0169f $ **FLOATING
C188 a_6092_17969.n23 VSS 0.0169f $ **FLOATING
C189 a_6092_17969.n24 VSS 0.27782f $ **FLOATING
C190 a_6092_17969.n25 VSS 0.01399f $ **FLOATING
C191 a_6092_17969.t16 VSS 0.10358f $ **FLOATING
C192 a_6092_17969.n26 VSS 0.22159f $ **FLOATING
C193 a_6092_17969.n28 VSS 0.26009f $ **FLOATING
C194 a_6092_17969.t13 VSS 0.10358f $ **FLOATING
C195 a_6092_17969.t10 VSS 0.10358f $ **FLOATING
C196 a_6092_17969.n29 VSS 0.41703f $ **FLOATING
C197 a_6092_17969.n30 VSS 0.9758f $ **FLOATING
C198 a_6092_17969.n31 VSS 0.0169f $ **FLOATING
C199 a_6092_17969.n32 VSS 0.01161f $ **FLOATING
C200 a_6092_17969.t15 VSS 0.10358f $ **FLOATING
C201 a_6092_17969.n40 VSS 0.01126f $ **FLOATING
C202 a_6092_17969.t9 VSS 0.0547f $ **FLOATING
C203 a_6092_17969.t7 VSS 1.03028f $ **FLOATING
C204 a_6092_17969.n41 VSS 1.97223f $ **FLOATING
C205 a_6092_17969.n43 VSS 0.0169f $ **FLOATING
C206 a_6092_17969.n45 VSS 0.0169f $ **FLOATING
C207 a_6092_17969.n47 VSS 0.0169f $ **FLOATING
C208 a_6092_17969.n49 VSS 0.0169f $ **FLOATING
C209 a_6092_17969.n51 VSS 0.0169f $ **FLOATING
C210 a_6092_17969.n53 VSS 0.0169f $ **FLOATING
C211 a_6092_17969.n54 VSS 0.0169f $ **FLOATING
C212 a_6092_17969.n55 VSS 0.27782f $ **FLOATING
C213 a_6092_17969.n56 VSS 0.01399f $ **FLOATING
C214 a_6092_17969.t8 VSS 0.10358f $ **FLOATING
C215 a_6092_17969.n57 VSS 0.22159f $ **FLOATING
C216 a_6092_17969.n59 VSS 0.13321f $ **FLOATING
C217 a_6092_17969.n60 VSS 0.92748f $ **FLOATING
C218 a_6092_17969.t12 VSS 0.10358f $ **FLOATING
C219 a_6092_17969.t4 VSS 0.10358f $ **FLOATING
C220 a_6092_17969.n61 VSS 0.42733f $ **FLOATING
C221 a_6092_17969.n62 VSS 1.43858f $ **FLOATING
C222 a_6092_17969.t17 VSS 0.10358f $ **FLOATING
C223 a_6092_17969.t14 VSS 0.10358f $ **FLOATING
C224 a_6092_17969.n63 VSS 0.42733f $ **FLOATING
C225 a_6092_17969.n64 VSS 1.24419f $ **FLOATING
C226 a_6092_17969.t2 VSS 0.0148f $ **FLOATING
C227 a_6092_17969.t1 VSS 0.0148f $ **FLOATING
C228 a_6092_17969.n65 VSS 0.03121f $ **FLOATING
C229 a_6092_17969.t27 VSS 0.06438f $ **FLOATING
C230 a_6092_17969.t35 VSS 0.0643f $ **FLOATING
C231 a_6092_17969.n66 VSS 0.11938f $ **FLOATING
C232 a_6092_17969.t20 VSS 0.0643f $ **FLOATING
C233 a_6092_17969.n67 VSS 0.05551f $ **FLOATING
C234 a_6092_17969.n68 VSS 0.14431f $ **FLOATING
C235 a_6092_17969.t29 VSS 0.0643f $ **FLOATING
C236 a_6092_17969.n69 VSS 0.05551f $ **FLOATING
C237 a_6092_17969.t28 VSS 0.0643f $ **FLOATING
C238 a_6092_17969.n70 VSS 0.0636f $ **FLOATING
C239 a_6092_17969.t18 VSS 0.0643f $ **FLOATING
C240 a_6092_17969.n71 VSS 0.0636f $ **FLOATING
C241 a_6092_17969.t26 VSS 0.0643f $ **FLOATING
C242 a_6092_17969.n72 VSS 0.0636f $ **FLOATING
C243 a_6092_17969.t30 VSS 0.0643f $ **FLOATING
C244 a_6092_17969.n73 VSS 0.0636f $ **FLOATING
C245 a_6092_17969.t19 VSS 0.0643f $ **FLOATING
C246 a_6092_17969.n74 VSS 0.30004f $ **FLOATING
C247 a_6092_17969.t11 VSS 0.24213f $ **FLOATING
C248 a_6092_17969.n75 VSS 4.17418f $ **FLOATING
C249 a_6092_17969.n76 VSS 1.82897f $ **FLOATING
C250 a_6092_17969.t33 VSS 0.0643f $ **FLOATING
C251 a_6092_17969.n77 VSS 0.20023f $ **FLOATING
C252 a_6092_17969.t22 VSS 0.0643f $ **FLOATING
C253 a_6092_17969.n78 VSS 0.0636f $ **FLOATING
C254 a_6092_17969.t31 VSS 0.0643f $ **FLOATING
C255 a_6092_17969.n79 VSS 0.0636f $ **FLOATING
C256 a_6092_17969.t34 VSS 0.0643f $ **FLOATING
C257 a_6092_17969.n80 VSS 0.0636f $ **FLOATING
C258 a_6092_17969.t24 VSS 0.0643f $ **FLOATING
C259 a_6092_17969.n81 VSS 0.0636f $ **FLOATING
C260 a_6092_17969.t23 VSS 0.0643f $ **FLOATING
C261 a_6092_17969.n82 VSS 0.05551f $ **FLOATING
C262 a_6092_17969.t25 VSS 0.06438f $ **FLOATING
C263 a_6092_17969.t21 VSS 0.0643f $ **FLOATING
C264 a_6092_17969.n83 VSS 0.11938f $ **FLOATING
C265 a_6092_17969.t32 VSS 0.0643f $ **FLOATING
C266 a_6092_17969.n84 VSS 0.05551f $ **FLOATING
C267 a_6092_17969.n85 VSS 0.14431f $ **FLOATING
C268 a_6092_17969.t0 VSS 0.0148f $ **FLOATING
C269 a_6092_17969.n86 VSS 0.03121f $ **FLOATING
C270 a_6092_17969.t3 VSS 0.0148f $ **FLOATING
C271 VDD.t62 VSS 0.02868f $ **FLOATING
C272 VDD.n0 VSS 0.01614f $ **FLOATING
C273 VDD.n1 VSS 0.1094f $ **FLOATING
C274 VDD.t60 VSS 0.03362f $ **FLOATING
C275 VDD.n2 VSS 0.08709f $ **FLOATING
C276 VDD.n3 VSS 0.01714f $ **FLOATING
C277 VDD.n4 VSS 0.18178f $ **FLOATING
C278 VDD.n5 VSS 0.01714f $ **FLOATING
C279 VDD.n6 VSS 0.12277f $ **FLOATING
C280 VDD.n7 VSS 0.01714f $ **FLOATING
C281 VDD.n8 VSS 0.12277f $ **FLOATING
C282 VDD.n9 VSS 0.01714f $ **FLOATING
C283 VDD.n10 VSS 0.16127f $ **FLOATING
C284 VDD.n11 VSS 0.05109f $ **FLOATING
C285 VDD.n12 VSS 0.01982f $ **FLOATING
C286 VDD.t45 VSS 0.02874f $ **FLOATING
C287 VDD.n13 VSS 0.07415f $ **FLOATING
C288 VDD.n14 VSS 0.02479f $ **FLOATING
C289 VDD.t40 VSS 0.03366f $ **FLOATING
C290 VDD.n15 VSS 0.019f $ **FLOATING
C291 VDD.n16 VSS 0.05818f $ **FLOATING
C292 VDD.t31 VSS 0.06597f $ **FLOATING
C293 VDD.n17 VSS 0.02436f $ **FLOATING
C294 VDD.n18 VSS 0.03986f $ **FLOATING
C295 VDD.t50 VSS 0.06595f $ **FLOATING
C296 VDD.n19 VSS 0.02479f $ **FLOATING
C297 VDD.n20 VSS 0.03986f $ **FLOATING
C298 VDD.t42 VSS 0.06599f $ **FLOATING
C299 VDD.n21 VSS 0.04395f $ **FLOATING
C300 VDD.n22 VSS 0.01982f $ **FLOATING
C301 VDD.n23 VSS 0.01612f $ **FLOATING
C302 VDD.t51 VSS 0.01547f $ **FLOATING
C303 VDD.n24 VSS 0.01612f $ **FLOATING
C304 VDD.t32 VSS 0.01547f $ **FLOATING
C305 VDD.n25 VSS 0.01614f $ **FLOATING
C306 VDD.t41 VSS 0.01547f $ **FLOATING
C307 VDD.n26 VSS 0.01614f $ **FLOATING
C308 VDD.n27 VSS 0.10538f $ **FLOATING
C309 VDD.n28 VSS 0.01714f $ **FLOATING
C310 VDD.n29 VSS 0.23646f $ **FLOATING
C311 VDD.n30 VSS 0.05109f $ **FLOATING
C312 VDD.t55 VSS 0.01547f $ **FLOATING
C313 VDD.n31 VSS 0.02436f $ **FLOATING
C314 VDD.n32 VSS 0.02479f $ **FLOATING
C315 VDD.t58 VSS 0.03366f $ **FLOATING
C316 VDD.t46 VSS 0.06599f $ **FLOATING
C317 VDD.t47 VSS 0.03647f $ **FLOATING
C318 VDD.n33 VSS 0.04395f $ **FLOATING
C319 VDD.n34 VSS 0.01612f $ **FLOATING
C320 VDD.n35 VSS 0.01982f $ **FLOATING
C321 VDD.n36 VSS 0.07415f $ **FLOATING
C322 VDD.n37 VSS 0.03986f $ **FLOATING
C323 VDD.t54 VSS 0.06595f $ **FLOATING
C324 VDD.n38 VSS 0.02479f $ **FLOATING
C325 VDD.n39 VSS 0.03986f $ **FLOATING
C326 VDD.t38 VSS 0.06597f $ **FLOATING
C327 VDD.n40 VSS 0.05818f $ **FLOATING
C328 VDD.n41 VSS 0.019f $ **FLOATING
C329 VDD.n42 VSS 0.01982f $ **FLOATING
C330 VDD.n43 VSS 0.01612f $ **FLOATING
C331 VDD.t39 VSS 0.01547f $ **FLOATING
C332 VDD.n44 VSS 0.01614f $ **FLOATING
C333 VDD.t59 VSS 0.01547f $ **FLOATING
C334 VDD.n45 VSS 0.01614f $ **FLOATING
C335 VDD.n46 VSS 0.0799f $ **FLOATING
C336 VDD.n47 VSS 0.07717f $ **FLOATING
C337 VDD.n51 VSS 0.64858f $ **FLOATING
C338 VDD.n65 VSS 0.01297f $ **FLOATING
C339 VDD.t29 VSS 0.1901f $ **FLOATING
C340 VDD.n68 VSS 0.35504f $ **FLOATING
C341 VDD.n69 VSS 0.51159f $ **FLOATING
C342 VDD.n70 VSS 0.01297f $ **FLOATING
C343 VDD.n82 VSS 0.01333f $ **FLOATING
C344 VDD.n83 VSS 0.01333f $ **FLOATING
C345 VDD.n84 VSS 0.01297f $ **FLOATING
C346 VDD.t34 VSS 0.1901f $ **FLOATING
C347 VDD.n90 VSS 0.36622f $ **FLOATING
C348 VDD.t22 VSS 0.1901f $ **FLOATING
C349 VDD.n97 VSS 0.3774f $ **FLOATING
C350 VDD.t0 VSS 0.1901f $ **FLOATING
C351 VDD.t14 VSS 0.1901f $ **FLOATING
C352 VDD.n107 VSS 0.3774f $ **FLOATING
C353 VDD.t5 VSS 0.1901f $ **FLOATING
C354 VDD.n114 VSS 0.36622f $ **FLOATING
C355 VDD.t2 VSS 0.1901f $ **FLOATING
C356 VDD.n119 VSS 0.01297f $ **FLOATING
C357 VDD.n120 VSS 0.01297f $ **FLOATING
C358 VDD.n121 VSS 0.35504f $ **FLOATING
C359 VDD.n123 VSS 0.01297f $ **FLOATING
C360 VDD.n135 VSS 0.01333f $ **FLOATING
C361 VDD.n164 VSS 0.01297f $ **FLOATING
C362 VDD.n165 VSS 0.01333f $ **FLOATING
C363 VDD.n212 VSS 0.01333f $ **FLOATING
C364 VDD.n213 VSS 0.01333f $ **FLOATING
C365 VDD.n215 VSS 0.64858f $ **FLOATING
C366 VDD.n216 VSS 0.51159f $ **FLOATING
C367 VDD.t43 VSS 0.1901f $ **FLOATING
C368 VDD.n217 VSS 0.22085f $ **FLOATING
C369 VDD.n223 VSS 0.21526f $ **FLOATING
C370 VDD.n224 VSS 0.36063f $ **FLOATING
C371 VDD.t7 VSS 0.1901f $ **FLOATING
C372 VDD.n225 VSS 0.20967f $ **FLOATING
C373 VDD.n231 VSS 0.20408f $ **FLOATING
C374 VDD.n232 VSS 0.37181f $ **FLOATING
C375 VDD.t11 VSS 0.1901f $ **FLOATING
C376 VDD.n233 VSS 0.19849f $ **FLOATING
C377 VDD.n239 VSS 0.19289f $ **FLOATING
C378 VDD.n240 VSS 0.3802f $ **FLOATING
C379 VDD.n241 VSS 0.19289f $ **FLOATING
C380 VDD.n247 VSS 0.19849f $ **FLOATING
C381 VDD.t17 VSS 0.1901f $ **FLOATING
C382 VDD.n248 VSS 0.37181f $ **FLOATING
C383 VDD.n249 VSS 0.20408f $ **FLOATING
C384 VDD.n255 VSS 0.20967f $ **FLOATING
C385 VDD.t3 VSS 0.1901f $ **FLOATING
C386 VDD.n256 VSS 0.36063f $ **FLOATING
C387 VDD.n257 VSS 0.21526f $ **FLOATING
C388 VDD.n263 VSS 0.22085f $ **FLOATING
C389 VDD.n266 VSS 0.01297f $ **FLOATING
C390 VDD.n267 VSS 0.01333f $ **FLOATING
C391 VDD.n268 VSS 0.01333f $ **FLOATING
C392 VDD.n303 VSS 0.02243f $ **FLOATING
C393 VDD.n304 VSS 0.13759f $ **FLOATING
C394 VDD.n305 VSS 0.05109f $ **FLOATING
C395 VDD.n306 VSS 0.01982f $ **FLOATING
C396 VDD.n307 VSS 0.04395f $ **FLOATING
C397 VDD.n308 VSS 0.02436f $ **FLOATING
C398 VDD.t65 VSS 0.02874f $ **FLOATING
C399 VDD.n309 VSS 0.03986f $ **FLOATING
C400 VDD.t56 VSS 0.03366f $ **FLOATING
C401 VDD.t48 VSS 0.06597f $ **FLOATING
C402 VDD.n310 VSS 0.05818f $ **FLOATING
C403 VDD.n311 VSS 0.019f $ **FLOATING
C404 VDD.n312 VSS 0.02479f $ **FLOATING
C405 VDD.t26 VSS 0.06595f $ **FLOATING
C406 VDD.n313 VSS 0.02479f $ **FLOATING
C407 VDD.t63 VSS 0.06599f $ **FLOATING
C408 VDD.n314 VSS 0.03986f $ **FLOATING
C409 VDD.n315 VSS 0.07415f $ **FLOATING
C410 VDD.n316 VSS 0.01982f $ **FLOATING
C411 VDD.n317 VSS 0.01612f $ **FLOATING
C412 VDD.t27 VSS 0.01547f $ **FLOATING
C413 VDD.n318 VSS 0.01612f $ **FLOATING
C414 VDD.t49 VSS 0.01547f $ **FLOATING
C415 VDD.n319 VSS 0.01614f $ **FLOATING
C416 VDD.t57 VSS 0.01547f $ **FLOATING
C417 VDD.n320 VSS 0.01614f $ **FLOATING
C418 VDD.n321 VSS 0.10554f $ **FLOATING
C419 VDD.n322 VSS 0.01714f $ **FLOATING
C420 VDD.n323 VSS 0.2372f $ **FLOATING
C421 VDD.n324 VSS 0.05109f $ **FLOATING
C422 VDD.t35 VSS 0.01547f $ **FLOATING
C423 VDD.n325 VSS 0.019f $ **FLOATING
C424 VDD.n326 VSS 0.07415f $ **FLOATING
C425 VDD.n327 VSS 0.03986f $ **FLOATING
C426 VDD.t66 VSS 0.06599f $ **FLOATING
C427 VDD.t67 VSS 0.03647f $ **FLOATING
C428 VDD.n328 VSS 0.01612f $ **FLOATING
C429 VDD.n329 VSS 0.01982f $ **FLOATING
C430 VDD.n330 VSS 0.04395f $ **FLOATING
C431 VDD.n331 VSS 0.02479f $ **FLOATING
C432 VDD.t33 VSS 0.06595f $ **FLOATING
C433 VDD.n332 VSS 0.02479f $ **FLOATING
C434 VDD.t36 VSS 0.03366f $ **FLOATING
C435 VDD.n333 VSS 0.05818f $ **FLOATING
C436 VDD.t52 VSS 0.06597f $ **FLOATING
C437 VDD.n334 VSS 0.03986f $ **FLOATING
C438 VDD.n335 VSS 0.02436f $ **FLOATING
C439 VDD.n336 VSS 0.01982f $ **FLOATING
C440 VDD.n337 VSS 0.01612f $ **FLOATING
C441 VDD.t53 VSS 0.01547f $ **FLOATING
C442 VDD.n338 VSS 0.01614f $ **FLOATING
C443 VDD.t37 VSS 0.01547f $ **FLOATING
C444 VDD.n339 VSS 0.01614f $ **FLOATING
C445 VDD.n340 VSS 0.0799f $ **FLOATING
C446 VDD.n341 VSS 0.09688f $ **FLOATING
C447 VDD.n342 VSS 0.01771f $ **FLOATING
C448 VDD.n343 VSS 0.01714f $ **FLOATING
C449 VDD.n344 VSS 0.31324f $ **FLOATING
C450 VDD.n345 VSS 0.01714f $ **FLOATING
C451 VDD.n346 VSS 0.12277f $ **FLOATING
C452 VDD.n347 VSS 0.01714f $ **FLOATING
C453 VDD.n348 VSS 0.12277f $ **FLOATING
C454 VDD.t30 VSS 0.03641f $ **FLOATING
C455 VDD.t69 VSS 0.01265f $ **FLOATING
C456 VDD.n349 VSS 0.01131f $ **FLOATING
C457 VDD.t28 VSS 0.03362f $ **FLOATING
C458 VDD.n350 VSS 0.18166f $ **FLOATING
C459 VDD.n351 VSS 0.10029f $ **FLOATING
C460 VDD.n352 VSS 0.40357f $ **FLOATING
C461 VDD.n353 VSS 0.26328f $ **FLOATING
C462 VDD.n354 VSS 0.18047f $ **FLOATING
C463 a_6681_14134.t13 VSS 0.1489f $ **FLOATING
C464 a_6681_14134.t15 VSS 0.1489f $ **FLOATING
C465 a_6681_14134.n0 VSS 0.82638f $ **FLOATING
C466 a_6681_14134.t18 VSS 0.1489f $ **FLOATING
C467 a_6681_14134.t16 VSS 0.1489f $ **FLOATING
C468 a_6681_14134.n1 VSS 0.61428f $ **FLOATING
C469 a_6681_14134.n2 VSS 3.04468f $ **FLOATING
C470 a_6681_14134.n3 VSS 0.02429f $ **FLOATING
C471 a_6681_14134.n4 VSS 0.01669f $ **FLOATING
C472 a_6681_14134.t19 VSS 0.1489f $ **FLOATING
C473 a_6681_14134.n5 VSS 0.02011f $ **FLOATING
C474 a_6681_14134.t6 VSS 0.07864f $ **FLOATING
C475 a_6681_14134.t4 VSS 1.4811f $ **FLOATING
C476 a_6681_14134.n12 VSS 2.83522f $ **FLOATING
C477 a_6681_14134.n13 VSS 0.39939f $ **FLOATING
C478 a_6681_14134.n14 VSS 0.01619f $ **FLOATING
C479 a_6681_14134.n15 VSS 0.02429f $ **FLOATING
C480 a_6681_14134.n17 VSS 0.02429f $ **FLOATING
C481 a_6681_14134.n19 VSS 0.02429f $ **FLOATING
C482 a_6681_14134.n21 VSS 0.02429f $ **FLOATING
C483 a_6681_14134.n23 VSS 0.02429f $ **FLOATING
C484 a_6681_14134.n25 VSS 0.02429f $ **FLOATING
C485 a_6681_14134.n26 VSS 0.02429f $ **FLOATING
C486 a_6681_14134.t5 VSS 0.1489f $ **FLOATING
C487 a_6681_14134.n29 VSS 0.31856f $ **FLOATING
C488 a_6681_14134.n30 VSS 0.0105f $ **FLOATING
C489 a_6681_14134.n31 VSS 0.37397f $ **FLOATING
C490 a_6681_14134.t17 VSS 0.1489f $ **FLOATING
C491 a_6681_14134.t14 VSS 0.1489f $ **FLOATING
C492 a_6681_14134.n32 VSS 0.59955f $ **FLOATING
C493 a_6681_14134.n33 VSS 1.40267f $ **FLOATING
C494 a_6681_14134.n34 VSS 0.02429f $ **FLOATING
C495 a_6681_14134.n35 VSS 0.01669f $ **FLOATING
C496 a_6681_14134.t8 VSS 0.22754f $ **FLOATING
C497 a_6681_14134.n36 VSS 0.02011f $ **FLOATING
C498 a_6681_14134.t7 VSS 1.4811f $ **FLOATING
C499 a_6681_14134.n43 VSS 2.83522f $ **FLOATING
C500 a_6681_14134.n44 VSS 0.39939f $ **FLOATING
C501 a_6681_14134.n45 VSS 0.01619f $ **FLOATING
C502 a_6681_14134.n46 VSS 0.02429f $ **FLOATING
C503 a_6681_14134.n48 VSS 0.02429f $ **FLOATING
C504 a_6681_14134.n50 VSS 0.02429f $ **FLOATING
C505 a_6681_14134.n52 VSS 0.02429f $ **FLOATING
C506 a_6681_14134.n54 VSS 0.02429f $ **FLOATING
C507 a_6681_14134.n56 VSS 0.02429f $ **FLOATING
C508 a_6681_14134.n57 VSS 0.02429f $ **FLOATING
C509 a_6681_14134.t20 VSS 0.1489f $ **FLOATING
C510 a_6681_14134.n60 VSS 0.31856f $ **FLOATING
C511 a_6681_14134.n61 VSS 0.0105f $ **FLOATING
C512 a_6681_14134.n62 VSS 0.1915f $ **FLOATING
C513 a_6681_14134.n63 VSS 0.35551f $ **FLOATING
C514 a_6681_14134.n64 VSS 2.01156f $ **FLOATING
C515 a_6681_14134.t0 VSS 0.09244f $ **FLOATING
C516 a_6681_14134.t22 VSS 0.09244f $ **FLOATING
C517 a_6681_14134.n65 VSS 1.20245f $ **FLOATING
C518 a_6681_14134.t2 VSS 0.09244f $ **FLOATING
C519 a_6681_14134.t21 VSS 0.09244f $ **FLOATING
C520 a_6681_14134.t12 VSS 0.02127f $ **FLOATING
C521 a_6681_14134.t10 VSS 0.02127f $ **FLOATING
C522 a_6681_14134.n66 VSS 0.04453f $ **FLOATING
C523 a_6681_14134.t24 VSS 0.09244f $ **FLOATING
C524 a_6681_14134.t9 VSS 0.09244f $ **FLOATING
C525 a_6681_14134.n68 VSS 0.23445f $ **FLOATING
C526 a_6681_14134.t11 VSS 0.09244f $ **FLOATING
C527 a_6681_14134.n69 VSS 0.24462f $ **FLOATING
C528 a_6681_14134.t23 VSS 0.09244f $ **FLOATING
C529 a_6681_14134.n70 VSS 0.24462f $ **FLOATING
C530 a_6681_14134.n71 VSS 0.23445f $ **FLOATING
C531 a_6681_14134.t3 VSS 0.02127f $ **FLOATING
C532 a_6681_14134.n72 VSS 0.04453f $ **FLOATING
C533 a_6681_14134.t1 VSS 0.02127f $ **FLOATING
C534 a_6681_4767.t27 VSS 0.04421f $ **FLOATING
C535 a_6681_4767.t12 VSS 0.01895f $ **FLOATING
C536 a_6681_4767.t18 VSS 0.01895f $ **FLOATING
C537 a_6681_4767.n9 VSS 0.04475f $ **FLOATING
C538 a_6681_4767.n10 VSS 0.16025f $ **FLOATING
C539 a_6681_4767.t17 VSS 0.01895f $ **FLOATING
C540 a_6681_4767.t24 VSS 0.01895f $ **FLOATING
C541 a_6681_4767.n11 VSS 0.04475f $ **FLOATING
C542 a_6681_4767.t8 VSS 0.01895f $ **FLOATING
C543 a_6681_4767.t23 VSS 0.01895f $ **FLOATING
C544 a_6681_4767.n12 VSS 0.04475f $ **FLOATING
C545 a_6681_4767.t4 VSS 0.01895f $ **FLOATING
C546 a_6681_4767.t20 VSS 0.01895f $ **FLOATING
C547 a_6681_4767.n13 VSS 0.04373f $ **FLOATING
C548 a_6681_4767.t14 VSS 0.01895f $ **FLOATING
C549 a_6681_4767.t21 VSS 0.01895f $ **FLOATING
C550 a_6681_4767.n14 VSS 0.04373f $ **FLOATING
C551 a_6681_4767.t10 VSS 0.01895f $ **FLOATING
C552 a_6681_4767.t15 VSS 0.01895f $ **FLOATING
C553 a_6681_4767.n15 VSS 0.04373f $ **FLOATING
C554 a_6681_4767.t25 VSS 0.01895f $ **FLOATING
C555 a_6681_4767.t9 VSS 0.01895f $ **FLOATING
C556 a_6681_4767.n16 VSS 0.04373f $ **FLOATING
C557 a_6681_4767.t3 VSS 0.01895f $ **FLOATING
C558 a_6681_4767.t26 VSS 0.01895f $ **FLOATING
C559 a_6681_4767.n17 VSS 0.04373f $ **FLOATING
C560 a_6681_4767.t19 VSS 0.01895f $ **FLOATING
C561 a_6681_4767.t13 VSS 0.01895f $ **FLOATING
C562 a_6681_4767.n18 VSS 0.04373f $ **FLOATING
C563 a_6681_4767.t22 VSS 0.01895f $ **FLOATING
C564 a_6681_4767.t16 VSS 0.01895f $ **FLOATING
C565 a_6681_4767.n19 VSS 0.04475f $ **FLOATING
C566 a_6681_4767.t7 VSS 0.01895f $ **FLOATING
C567 a_6681_4767.t6 VSS 0.01895f $ **FLOATING
C568 a_6681_4767.n20 VSS 0.04475f $ **FLOATING
C569 a_6681_4767.t5 VSS 0.01895f $ **FLOATING
C570 a_6681_4767.t11 VSS 0.01895f $ **FLOATING
C571 a_6681_4767.n21 VSS 0.04475f $ **FLOATING
C572 a_6681_4767.n22 VSS 0.18025f $ **FLOATING
C573 a_6681_4767.n23 VSS 0.18025f $ **FLOATING
C574 a_6681_4767.n24 VSS 0.43966f $ **FLOATING
C575 a_6681_4767.n25 VSS 0.42532f $ **FLOATING
C576 a_6681_4767.n26 VSS 0.17285f $ **FLOATING
C577 a_6681_4767.n27 VSS 0.17285f $ **FLOATING
C578 a_6681_4767.n28 VSS 0.17285f $ **FLOATING
C579 a_6681_4767.n29 VSS 0.17285f $ **FLOATING
C580 a_6681_4767.n30 VSS 0.44215f $ **FLOATING
C581 a_6681_4767.n31 VSS 0.44955f $ **FLOATING
C582 a_6681_4767.n32 VSS 0.16879f $ **FLOATING
C583 a_6681_4767.n33 VSS 0.04604f $ **FLOATING
C584 a_6681_4767.n34 VSS 0.02203f $ **FLOATING
C585 a_6681_4767.t1 VSS 0.04421f $ **FLOATING
C586 a_6681_4767.n48 VSS 0.09459f $ **FLOATING
C587 a_6681_4767.n52 VSS 0.11859f $ **FLOATING
C588 a_6681_4767.t0 VSS 0.4397f $ **FLOATING
C589 a_6681_4767.n53 VSS 0.70858f $ **FLOATING
C590 a_6681_4767.n54 VSS 0.12689f $ **FLOATING
C591 a_6681_4767.t2 VSS 0.02158f $ **FLOATING
C592 a_4943_7756.t7 VSS 0.02923f $ **FLOATING
C593 a_4943_7756.t31 VSS 0.21262f $ **FLOATING
C594 a_4943_7756.t14 VSS 0.21141f $ **FLOATING
C595 a_4943_7756.t26 VSS 0.21132f $ **FLOATING
C596 a_4943_7756.n9 VSS 0.11994f $ **FLOATING
C597 a_4943_7756.n10 VSS 0.14799f $ **FLOATING
C598 a_4943_7756.t25 VSS 0.21141f $ **FLOATING
C599 a_4943_7756.t35 VSS 0.21132f $ **FLOATING
C600 a_4943_7756.n11 VSS 0.11994f $ **FLOATING
C601 a_4943_7756.n12 VSS 0.02095f $ **FLOATING
C602 a_4943_7756.t39 VSS 0.21141f $ **FLOATING
C603 a_4943_7756.t13 VSS 0.21132f $ **FLOATING
C604 a_4943_7756.n13 VSS 0.11994f $ **FLOATING
C605 a_4943_7756.n14 VSS 0.02095f $ **FLOATING
C606 a_4943_7756.t40 VSS 0.21141f $ **FLOATING
C607 a_4943_7756.t15 VSS 0.21132f $ **FLOATING
C608 a_4943_7756.n15 VSS 0.11994f $ **FLOATING
C609 a_4943_7756.n16 VSS 0.02095f $ **FLOATING
C610 a_4943_7756.t41 VSS 0.21141f $ **FLOATING
C611 a_4943_7756.t17 VSS 0.21132f $ **FLOATING
C612 a_4943_7756.n17 VSS 0.11994f $ **FLOATING
C613 a_4943_7756.n18 VSS 0.02095f $ **FLOATING
C614 a_4943_7756.n19 VSS 0.02095f $ **FLOATING
C615 a_4943_7756.t30 VSS 0.21141f $ **FLOATING
C616 a_4943_7756.n20 VSS 0.0113f $ **FLOATING
C617 a_4943_7756.t33 VSS 0.21141f $ **FLOATING
C618 a_4943_7756.n21 VSS 0.07214f $ **FLOATING
C619 a_4943_7756.n22 VSS 0.04736f $ **FLOATING
C620 a_4943_7756.t3 VSS 0.16079f $ **FLOATING
C621 a_4943_7756.t4 VSS 0.01253f $ **FLOATING
C622 a_4943_7756.t6 VSS 0.01253f $ **FLOATING
C623 a_4943_7756.n42 VSS 0.02505f $ **FLOATING
C624 a_4943_7756.n45 VSS 0.1113f $ **FLOATING
C625 a_4943_7756.t5 VSS 0.16079f $ **FLOATING
C626 a_4943_7756.n46 VSS 0.04736f $ **FLOATING
C627 a_4943_7756.n47 VSS 0.07214f $ **FLOATING
C628 a_4943_7756.n48 VSS 0.02095f $ **FLOATING
C629 a_4943_7756.t22 VSS 0.21141f $ **FLOATING
C630 a_4943_7756.t32 VSS 0.21132f $ **FLOATING
C631 a_4943_7756.n49 VSS 0.11994f $ **FLOATING
C632 a_4943_7756.n50 VSS 0.02095f $ **FLOATING
C633 a_4943_7756.t23 VSS 0.21141f $ **FLOATING
C634 a_4943_7756.t34 VSS 0.21132f $ **FLOATING
C635 a_4943_7756.n51 VSS 0.11994f $ **FLOATING
C636 a_4943_7756.n52 VSS 0.02095f $ **FLOATING
C637 a_4943_7756.t10 VSS 0.21141f $ **FLOATING
C638 a_4943_7756.t21 VSS 0.21132f $ **FLOATING
C639 a_4943_7756.n53 VSS 0.11994f $ **FLOATING
C640 a_4943_7756.n54 VSS 0.02095f $ **FLOATING
C641 a_4943_7756.t38 VSS 0.21141f $ **FLOATING
C642 a_4943_7756.t12 VSS 0.21132f $ **FLOATING
C643 a_4943_7756.n55 VSS 0.11994f $ **FLOATING
C644 a_4943_7756.n56 VSS 0.02095f $ **FLOATING
C645 a_4943_7756.t11 VSS 0.21141f $ **FLOATING
C646 a_4943_7756.t24 VSS 0.21132f $ **FLOATING
C647 a_4943_7756.n57 VSS 0.11994f $ **FLOATING
C648 a_4943_7756.n58 VSS 0.02095f $ **FLOATING
C649 a_4943_7756.t18 VSS 0.21218f $ **FLOATING
C650 a_4943_7756.n59 VSS 0.12882f $ **FLOATING
C651 a_4943_7756.t20 VSS 0.2127f $ **FLOATING
C652 a_4943_7756.t29 VSS 0.21218f $ **FLOATING
C653 a_4943_7756.n60 VSS 0.23123f $ **FLOATING
C654 a_4943_7756.t43 VSS 0.21218f $ **FLOATING
C655 a_4943_7756.n61 VSS 0.08346f $ **FLOATING
C656 a_4943_7756.t8 VSS 0.21218f $ **FLOATING
C657 a_4943_7756.n62 VSS 0.08346f $ **FLOATING
C658 a_4943_7756.t9 VSS 0.21218f $ **FLOATING
C659 a_4943_7756.n63 VSS 0.08346f $ **FLOATING
C660 a_4943_7756.t37 VSS 0.21218f $ **FLOATING
C661 a_4943_7756.n64 VSS 0.08346f $ **FLOATING
C662 a_4943_7756.t36 VSS 0.21218f $ **FLOATING
C663 a_4943_7756.n65 VSS 0.08346f $ **FLOATING
C664 a_4943_7756.t27 VSS 0.21218f $ **FLOATING
C665 a_4943_7756.n66 VSS 0.08346f $ **FLOATING
C666 a_4943_7756.t28 VSS 0.21218f $ **FLOATING
C667 a_4943_7756.n67 VSS 0.08346f $ **FLOATING
C668 a_4943_7756.t16 VSS 0.21218f $ **FLOATING
C669 a_4943_7756.n68 VSS 0.08346f $ **FLOATING
C670 a_4943_7756.t42 VSS 0.21218f $ **FLOATING
C671 a_4943_7756.n69 VSS 0.08346f $ **FLOATING
C672 a_4943_7756.t19 VSS 0.21218f $ **FLOATING
C673 a_4943_7756.n70 VSS 0.14747f $ **FLOATING
C674 a_4943_7756.n71 VSS 0.24566f $ **FLOATING
C675 a_4943_7756.n72 VSS 0.06486f $ **FLOATING
C676 a_4943_7756.t1 VSS 0.02923f $ **FLOATING
C677 a_4943_7756.n86 VSS 0.06253f $ **FLOATING
C678 a_4943_7756.n90 VSS 0.0784f $ **FLOATING
C679 a_4943_7756.t0 VSS 0.29068f $ **FLOATING
C680 a_4943_7756.n91 VSS 0.46844f $ **FLOATING
C681 a_4943_7756.n92 VSS 0.08389f $ **FLOATING
C682 a_4943_7756.t2 VSS 0.01427f $ **FLOATING
.ends
