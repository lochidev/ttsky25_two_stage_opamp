* NGSPICE file created from two_stage_op_amp.ext - technology: sky130A

.subckt two_stage_op_amp IBIAS EN VOUT VDD VN VP VSS
X0 VSS.t104 VSS.t103 VSS.t104 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X1 VDD.t71 a_2479_7336.t18 VOUT.t16 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X2 VSS.t132 a_2080_2896.t6 a_2080_2896.t7 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X3 VDD.t70 a_2479_7336.t19 VOUT.t12 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X4 VDD.t52 VDD.t51 VDD.t52 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X5 VSS.t124 a_2080_2896.t8 a_4920_2896.t23 VSS.t107 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 VSS.t115 a_2080_2896.t9 a_4920_2896.t22 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X7 a_2479_7336.t8 a_2479_7336.t7 a_2479_7336.t8 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X8 VSS.t102 VSS.t101 VSS.t102 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X9 VDD.t50 VDD.t49 VDD.t50 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X10 VDD.t69 a_2479_7336.t20 VOUT.t14 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X11 VDD.t68 a_2479_7336.t21 VOUT.t6 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X12 a_4920_2896.t21 a_2080_2896.t10 VSS.t138 VSS.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X13 a_2479_7336.t6 a_2479_7336.t4 a_2479_7336.t5 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X14 a_2479_7336.t12 VP.t0 a_2995_7336.t8 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X15 VSS.t22 a_2080_2896.t11 a_4920_2896.t20 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 VSS.t100 VSS.t99 VSS.t100 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X17 a_2995_7336.t13 VN.t0 a_2479_9004.t20 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X18 VDD.t67 a_2479_7336.t22 VOUT.t2 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X19 a_2479_9004.t19 VN.t1 a_2995_7336.t10 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X20 VSS.t98 VSS.t97 VSS.t98 VSS.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X21 a_2479_9004.t4 a_2479_9004.t3 a_2479_9004.t4 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X22 VSS.t96 VSS.t95 VSS.t96 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X23 a_4920_2896.t19 a_2080_2896.t12 VSS.t32 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X24 a_2479_9004.t2 a_2479_9004.t0 a_2479_9004.t1 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X25 a_2479_9004.t18 VN.t2 a_2995_7336.t16 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X26 VSS.t133 a_2080_2896.t13 a_4920_2896.t18 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X27 VOUT.t1 a_2479_7336.t23 VDD.t66 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X28 VSS.t94 VSS.t93 VSS.t94 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X29 VDD.t48 VDD.t46 VDD.t48 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X30 a_2995_7336.t7 VP.t1 a_2479_7336.t2 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X31 VSS.t92 VSS.t91 VSS.t92 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X32 a_3758_2896.t11 a_2080_2896.t14 VSS.t135 VSS.t107 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X33 a_4920_2896.t17 a_2080_2896.t15 VSS.t137 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X34 a_2479_7336.t1 VP.t2 a_2995_7336.t6 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X35 a_3758_2896.t10 a_2080_2896.t16 VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X36 VOUT.t11 a_2479_7336.t24 VDD.t65 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X37 VSS.t131 a_2080_2896.t17 a_3758_2896.t9 VSS.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X38 a_4920_2896.t26 a_4920_2896.t25 a_4920_2896.t26 VSS.t127 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X39 a_4920_2896.t16 a_2080_2896.t18 VSS.t4 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X40 a_3758_2896.t8 a_2080_2896.t19 VSS.t8 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X41 a_3758_2896.t7 a_2080_2896.t20 VSS.t109 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X42 a_4920_2896.t24 EN.t0 VOUT.t0 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X43 a_2995_7336.t5 VP.t3 a_2479_7336.t10 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X44 VDD.t72 a_2479_9004.t11 a_2479_9004.t12 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X45 VOUT.t31 VOUT.t29 VOUT.t30 VSS.t116 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X46 a_4920_2896.t15 a_2080_2896.t21 VSS.t111 VSS.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X47 VDD.t45 VDD.t44 VDD.t45 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X48 VSS.t123 a_2080_2896.t22 a_4920_2896.t14 VSS.t120 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X49 VDD.t43 VDD.t42 VDD.t43 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X50 VSS.t90 VSS.t89 VSS.t90 VSS.t79 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X51 VDD.t64 a_2479_7336.t25 VOUT.t3 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X52 VSS.t88 VSS.t86 VSS.t87 VSS.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X53 VSS.t85 VSS.t84 VSS.t85 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X54 VOUT.t28 VOUT.t26 VOUT.t27 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X55 VSS.t114 a_2080_2896.t23 a_4920_2896.t13 VSS.t113 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X56 VOUT.t25 VOUT.t24 VOUT.t25 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X57 a_2995_7336.t0 VN.t3 a_2479_9004.t17 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X58 VDD.t63 a_2479_7336.t26 VOUT.t13 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X59 VSS.t83 VSS.t81 VSS.t82 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X60 VDD.t41 VDD.t39 VDD.t40 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X61 a_2479_9004.t10 a_2479_9004.t9 VDD.t73 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X62 mim_cap_0.C1.t1 VOUT.t19 sky130_fd_pr__cap_mim_m3_1 l=25.5 w=25.5
X63 VDD.t62 a_2479_7336.t27 VOUT.t4 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X64 VSS.t7 a_2080_2896.t24 a_3758_2896.t6 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X65 a_4920_2896.t12 a_2080_2896.t25 VSS.t1 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X66 VSS.t80 VSS.t78 VSS.t80 VSS.t79 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X67 VOUT.t5 a_2479_7336.t28 VDD.t61 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X68 VDD.t76 a_2479_9004.t21 a_2479_7336.t15 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X69 VDD.t38 VDD.t37 VDD.t38 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X70 VSS.t77 VSS.t76 VSS.t77 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X71 VDD.t36 VDD.t35 VDD.t36 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X72 VOUT.t9 a_2479_7336.t29 VDD.t60 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X73 VSS.t122 a_2080_2896.t26 a_3758_2896.t5 VSS.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X74 VSS.t75 VSS.t74 VSS.t75 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X75 VDD.t34 VDD.t33 VDD.t34 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X76 VSS.t73 VSS.t72 VSS.t73 VSS.t51 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X77 VDD.t32 VDD.t30 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X78 a_3758_2896.t4 a_2080_2896.t27 VSS.t121 VSS.t120 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X79 VSS.t71 VSS.t70 VSS.t71 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X80 VSS.t69 VSS.t68 VSS.t69 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X81 VSS.t67 VSS.t66 VSS.t67 VSS.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X82 a_2995_7336.t4 VP.t4 a_2479_7336.t9 VSS.t79 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X83 VSS.t65 VSS.t64 VSS.t65 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X84 a_4920_2896.t11 a_2080_2896.t28 VSS.t119 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X85 a_2479_7336.t16 VP.t5 a_2995_7336.t3 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X86 a_2080_2896.t3 a_2080_2896.t1 a_2080_2896.t2 VSS.t112 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X87 a_2479_7336.t3 a_2479_9004.t22 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X88 VSS.t118 a_2080_2896.t29 a_4920_2896.t10 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X89 a_2995_7336.t15 VN.t4 a_2479_9004.t16 VSS.t51 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X90 VOUT.t8 a_2479_7336.t30 VDD.t59 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X91 a_4920_2896.t9 a_2080_2896.t30 VSS.t117 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X92 a_2479_9004.t15 VN.t5 a_2995_7336.t11 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X93 VDD.t74 a_2479_9004.t23 a_2479_7336.t13 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X94 VDD.t29 VDD.t27 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X95 VSS.t108 a_2080_2896.t31 a_4920_2896.t8 VSS.t107 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X96 VOUT.t18 a_2479_7336.t31 VDD.t58 VDD.t47 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X97 VSS.t106 a_2080_2896.t32 a_4920_2896.t7 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X98 a_2995_7336.t12 VN.t6 a_2479_9004.t14 VSS.t79 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X99 VDD.t26 VDD.t24 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X100 a_4920_2896.t6 a_2080_2896.t33 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X101 a_2479_9004.t13 VN.t7 a_2995_7336.t9 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X102 VSS.t6 a_2080_2896.t34 a_4920_2896.t5 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X103 VSS.t63 VSS.t61 VSS.t63 VSS.t62 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X104 a_2995_7336.t2 VP.t6 a_2479_7336.t11 VSS.t51 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X105 a_2479_7336.t0 VP.t7 a_2995_7336.t1 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X106 VSS.t60 VSS.t58 VSS.t60 VSS.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X107 VSS.t21 a_2080_2896.t35 a_3758_2896.t3 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X108 VSS.t134 a_2080_2896.t36 a_3758_2896.t2 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X109 VSS.t57 VSS.t55 VSS.t56 VSS.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X110 a_3758_2896.t1 a_2080_2896.t37 VSS.t16 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X111 VDD.t1 a_2479_9004.t7 a_2479_9004.t8 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X112 VSS.t24 a_2080_2896.t38 a_3758_2896.t0 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X113 IBIAS.t2 IBIAS.t1 IBIAS.t2 VSS.t129 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X114 VSS.t54 VSS.t53 VSS.t54 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X115 VDD.t23 VDD.t22 VDD.t23 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X116 VSS.t130 a_2080_2896.t39 a_4920_2896.t4 VSS.t113 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X117 VDD.t21 VDD.t19 VDD.t20 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X118 IBIAS.t0 EN.t1 a_2080_2896.t0 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X119 VSS.t52 VSS.t50 VSS.t52 VSS.t51 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X120 a_2479_7336.t14 a_2479_9004.t24 VDD.t75 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X121 a_4920_2896.t3 a_2080_2896.t40 VSS.t27 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X122 a_4920_2896.t2 a_2080_2896.t41 VSS.t105 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X123 VOUT.t7 a_2479_7336.t32 VDD.t57 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X124 a_2479_7336.t17 mim_cap_0.C1.t0 VSS.t128 sky130_fd_pr__res_xhigh_po_1p41 l=14
X125 VDD.t18 VDD.t16 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X126 VDD.t15 VDD.t13 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X127 a_3758_2896.t13 a_3758_2896.t12 a_3758_2896.t13 VSS.t126 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X128 VOUT.t15 a_2479_7336.t33 VDD.t56 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X129 VOUT.t23 VOUT.t22 VOUT.t23 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X130 a_4920_2896.t1 a_2080_2896.t42 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X131 a_3758_2896.t14 EN.t2 a_2995_7336.t14 VSS.t110 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X132 VSS.t125 a_2080_2896.t43 a_4920_2896.t0 VSS.t120 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X133 VOUT.t21 VOUT.t20 VOUT.t21 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X134 VOUT.t17 a_2479_7336.t34 VDD.t54 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X135 VSS.t49 VSS.t46 VSS.t48 VSS.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X136 a_2995_7336.t19 a_2995_7336.t17 a_2995_7336.t18 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X137 VDD.t12 VDD.t10 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X138 VSS.t45 VSS.t44 VSS.t45 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X139 VDD.t9 VDD.t6 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X140 a_2080_2896.t5 a_2080_2896.t4 VSS.t136 VSS.t113 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X141 VSS.t43 VSS.t41 VSS.t42 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X142 VSS.t40 VSS.t38 VSS.t40 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X143 VDD.t53 a_2479_7336.t35 VOUT.t10 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X144 VSS.t37 VSS.t35 VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X145 a_2479_9004.t6 a_2479_9004.t5 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X146 VSS.t34 VSS.t33 VSS.t34 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
C0 VP VN 5.95617f
C1 EN IBIAS 0.80152f
C2 VDD VOUT 9.55719f
C3 VOUT VN 0.15325f
C4 EN VOUT 0.69581f
C5 VDD mim_cap_0.C1 0.11752f
C6 VOUT mim_cap_0.C1 57.8517f
C7 VP VOUT 0.38099f
R0 VSS.n2095 VSS.n2094 2542.66
R1 VSS.n553 VSS.n538 1321.06
R2 VSS.n551 VSS.n540 1321.06
R3 VSS.n2096 VSS.n517 1321.06
R4 VSS.n634 VSS.n523 1321.06
R5 VSS.n1736 VSS.n876 1268.91
R6 VSS.n1817 VSS.n856 1268.91
R7 VSS.n1692 VSS.n1691 1268.91
R8 VSS.n1770 VSS.n854 1268.91
R9 VSS.n1449 VSS.n1393 1268.91
R10 VSS.n1538 VSS.n1119 1268.91
R11 VSS.n1411 VSS.n1149 1268.91
R12 VSS.n1495 VSS.n1494 1268.91
R13 VSS.n1557 VSS.n1049 1268.91
R14 VSS.n1665 VSS.n901 1268.91
R15 VSS.n1622 VSS.n1621 1268.91
R16 VSS.n1559 VSS.n1046 1268.91
R17 VSS.n424 VSS.n219 1182
R18 VSS.n2448 VSS.n101 1182
R19 VSS.n422 VSS.n221 1182
R20 VSS.n2392 VSS.n106 1182
R21 VSS.n2092 VSS.n647 1182
R22 VSS.n2017 VSS.n788 1182
R23 VSS.n1391 VSS.n1152 1182
R24 VSS.n1830 VSS.n838 1182
R25 VSS.n1973 VSS.n842 996.588
R26 VSS.n2095 VSS.n516 614.067
R27 VSS.n1925 VSS.n1924 602.588
R28 VSS.n1877 VSS.n1876 602.588
R29 VSS.n600 VSS.n599 585
R30 VSS.n599 VSS.n472 585
R31 VSS.n598 VSS.n471 585
R32 VSS.n2157 VSS.n471 585
R33 VSS.n597 VSS.n596 585
R34 VSS.n596 VSS.n467 585
R35 VSS.n595 VSS.n466 585
R36 VSS.n2163 VSS.n466 585
R37 VSS.n594 VSS.n465 585
R38 VSS.n2164 VSS.n465 585
R39 VSS.n593 VSS.n464 585
R40 VSS.n2165 VSS.n464 585
R41 VSS.n592 VSS.n591 585
R42 VSS.n591 VSS.n460 585
R43 VSS.n590 VSS.n459 585
R44 VSS.n2171 VSS.n459 585
R45 VSS.n589 VSS.n458 585
R46 VSS.n2172 VSS.n458 585
R47 VSS.n588 VSS.n457 585
R48 VSS.n2173 VSS.n457 585
R49 VSS.n587 VSS.n586 585
R50 VSS.n586 VSS.n453 585
R51 VSS.n585 VSS.n452 585
R52 VSS.n2179 VSS.n452 585
R53 VSS.n584 VSS.n451 585
R54 VSS.n2180 VSS.n451 585
R55 VSS.n583 VSS.n450 585
R56 VSS.n2181 VSS.n450 585
R57 VSS.n582 VSS.n581 585
R58 VSS.n581 VSS.n446 585
R59 VSS.n580 VSS.n445 585
R60 VSS.n2187 VSS.n445 585
R61 VSS.n579 VSS.n444 585
R62 VSS.n2188 VSS.n444 585
R63 VSS.n578 VSS.n443 585
R64 VSS.n2189 VSS.n443 585
R65 VSS.n577 VSS.n576 585
R66 VSS.n576 VSS.n437 585
R67 VSS.n575 VSS.n436 585
R68 VSS.n2195 VSS.n436 585
R69 VSS.n574 VSS.n573 585
R70 VSS.n573 VSS.n435 585
R71 VSS.n572 VSS.n525 585
R72 VSS.n572 VSS.n571 585
R73 VSS.n562 VSS.n526 585
R74 VSS.n527 VSS.n526 585
R75 VSS.n564 VSS.n563 585
R76 VSS.n565 VSS.n564 585
R77 VSS.n561 VSS.n532 585
R78 VSS.n532 VSS.n531 585
R79 VSS.n560 VSS.n559 585
R80 VSS.n559 VSS.n558 585
R81 VSS.n534 VSS.n533 585
R82 VSS.n535 VSS.n534 585
R83 VSS.n551 VSS.n550 585
R84 VSS.n552 VSS.n551 585
R85 VSS.n549 VSS.n540 585
R86 VSS.n548 VSS.n547 585
R87 VSS.n545 VSS.n541 585
R88 VSS.n543 VSS.n542 585
R89 VSS.n538 VSS.n537 585
R90 VSS.n539 VSS.n538 585
R91 VSS.n554 VSS.n553 585
R92 VSS.n553 VSS.n552 585
R93 VSS.n555 VSS.n536 585
R94 VSS.n536 VSS.n535 585
R95 VSS.n557 VSS.n556 585
R96 VSS.n558 VSS.n557 585
R97 VSS.n530 VSS.n529 585
R98 VSS.n531 VSS.n530 585
R99 VSS.n567 VSS.n566 585
R100 VSS.n566 VSS.n565 585
R101 VSS.n568 VSS.n528 585
R102 VSS.n528 VSS.n527 585
R103 VSS.n570 VSS.n569 585
R104 VSS.n571 VSS.n570 585
R105 VSS.n440 VSS.n438 585
R106 VSS.n438 VSS.n435 585
R107 VSS.n2194 VSS.n2193 585
R108 VSS.n2195 VSS.n2194 585
R109 VSS.n2192 VSS.n439 585
R110 VSS.n439 VSS.n437 585
R111 VSS.n2191 VSS.n2190 585
R112 VSS.n2190 VSS.n2189 585
R113 VSS.n442 VSS.n441 585
R114 VSS.n2188 VSS.n442 585
R115 VSS.n2186 VSS.n2185 585
R116 VSS.n2187 VSS.n2186 585
R117 VSS.n2184 VSS.n447 585
R118 VSS.n447 VSS.n446 585
R119 VSS.n2183 VSS.n2182 585
R120 VSS.n2182 VSS.n2181 585
R121 VSS.n449 VSS.n448 585
R122 VSS.n2180 VSS.n449 585
R123 VSS.n2178 VSS.n2177 585
R124 VSS.n2179 VSS.n2178 585
R125 VSS.n2176 VSS.n454 585
R126 VSS.n454 VSS.n453 585
R127 VSS.n2175 VSS.n2174 585
R128 VSS.n2174 VSS.n2173 585
R129 VSS.n456 VSS.n455 585
R130 VSS.n2172 VSS.n456 585
R131 VSS.n2170 VSS.n2169 585
R132 VSS.n2171 VSS.n2170 585
R133 VSS.n2168 VSS.n461 585
R134 VSS.n461 VSS.n460 585
R135 VSS.n2167 VSS.n2166 585
R136 VSS.n2166 VSS.n2165 585
R137 VSS.n463 VSS.n462 585
R138 VSS.n2164 VSS.n463 585
R139 VSS.n2162 VSS.n2161 585
R140 VSS.n2163 VSS.n2162 585
R141 VSS.n2160 VSS.n468 585
R142 VSS.n468 VSS.n467 585
R143 VSS.n2159 VSS.n2158 585
R144 VSS.n2158 VSS.n2157 585
R145 VSS.n470 VSS.n469 585
R146 VSS.n472 VSS.n470 585
R147 VSS.n2096 VSS.n518 585
R148 VSS.n2099 VSS.n2098 585
R149 VSS.n521 VSS.n520 585
R150 VSS.n2095 VSS.n521 585
R151 VSS.n524 VSS.n522 585
R152 VSS.n634 VSS.n633 585
R153 VSS.n632 VSS.n523 585
R154 VSS.n523 VSS.n516 585
R155 VSS.n631 VSS.n515 585
R156 VSS.n2107 VSS.n515 585
R157 VSS.n630 VSS.n514 585
R158 VSS.n2108 VSS.n514 585
R159 VSS.n629 VSS.n513 585
R160 VSS.n2109 VSS.n513 585
R161 VSS.n628 VSS.n627 585
R162 VSS.n627 VSS.n509 585
R163 VSS.n626 VSS.n508 585
R164 VSS.n2115 VSS.n508 585
R165 VSS.n625 VSS.n507 585
R166 VSS.n2116 VSS.n507 585
R167 VSS.n624 VSS.n506 585
R168 VSS.n2117 VSS.n506 585
R169 VSS.n623 VSS.n622 585
R170 VSS.n622 VSS.n502 585
R171 VSS.n621 VSS.n501 585
R172 VSS.n2123 VSS.n501 585
R173 VSS.n620 VSS.n500 585
R174 VSS.n2124 VSS.n500 585
R175 VSS.n619 VSS.n499 585
R176 VSS.n2125 VSS.n499 585
R177 VSS.n618 VSS.n617 585
R178 VSS.n617 VSS.n495 585
R179 VSS.n616 VSS.n494 585
R180 VSS.n2131 VSS.n494 585
R181 VSS.n615 VSS.n493 585
R182 VSS.n2132 VSS.n493 585
R183 VSS.n614 VSS.n492 585
R184 VSS.n2133 VSS.n492 585
R185 VSS.n613 VSS.n612 585
R186 VSS.n612 VSS.n488 585
R187 VSS.n611 VSS.n487 585
R188 VSS.n2139 VSS.n487 585
R189 VSS.n610 VSS.n486 585
R190 VSS.n2140 VSS.n486 585
R191 VSS.n609 VSS.n485 585
R192 VSS.n2141 VSS.n485 585
R193 VSS.n608 VSS.n607 585
R194 VSS.n607 VSS.n481 585
R195 VSS.n606 VSS.n480 585
R196 VSS.n2147 VSS.n480 585
R197 VSS.n605 VSS.n479 585
R198 VSS.n2148 VSS.n479 585
R199 VSS.n604 VSS.n478 585
R200 VSS.n2149 VSS.n478 585
R201 VSS.n603 VSS.n602 585
R202 VSS.n602 VSS.n474 585
R203 VSS.n601 VSS.n473 585
R204 VSS.n2155 VSS.n473 585
R205 VSS.n2154 VSS.n2153 585
R206 VSS.n2155 VSS.n2154 585
R207 VSS.n2152 VSS.n475 585
R208 VSS.n475 VSS.n474 585
R209 VSS.n2151 VSS.n2150 585
R210 VSS.n2150 VSS.n2149 585
R211 VSS.n477 VSS.n476 585
R212 VSS.n2148 VSS.n477 585
R213 VSS.n2146 VSS.n2145 585
R214 VSS.n2147 VSS.n2146 585
R215 VSS.n2144 VSS.n482 585
R216 VSS.n482 VSS.n481 585
R217 VSS.n2143 VSS.n2142 585
R218 VSS.n2142 VSS.n2141 585
R219 VSS.n484 VSS.n483 585
R220 VSS.n2140 VSS.n484 585
R221 VSS.n2138 VSS.n2137 585
R222 VSS.n2139 VSS.n2138 585
R223 VSS.n2136 VSS.n489 585
R224 VSS.n489 VSS.n488 585
R225 VSS.n2135 VSS.n2134 585
R226 VSS.n2134 VSS.n2133 585
R227 VSS.n491 VSS.n490 585
R228 VSS.n2132 VSS.n491 585
R229 VSS.n2130 VSS.n2129 585
R230 VSS.n2131 VSS.n2130 585
R231 VSS.n2128 VSS.n496 585
R232 VSS.n496 VSS.n495 585
R233 VSS.n2127 VSS.n2126 585
R234 VSS.n2126 VSS.n2125 585
R235 VSS.n498 VSS.n497 585
R236 VSS.n2124 VSS.n498 585
R237 VSS.n2122 VSS.n2121 585
R238 VSS.n2123 VSS.n2122 585
R239 VSS.n2120 VSS.n503 585
R240 VSS.n503 VSS.n502 585
R241 VSS.n2119 VSS.n2118 585
R242 VSS.n2118 VSS.n2117 585
R243 VSS.n505 VSS.n504 585
R244 VSS.n2116 VSS.n505 585
R245 VSS.n2114 VSS.n2113 585
R246 VSS.n2115 VSS.n2114 585
R247 VSS.n2112 VSS.n510 585
R248 VSS.n510 VSS.n509 585
R249 VSS.n2111 VSS.n2110 585
R250 VSS.n2110 VSS.n2109 585
R251 VSS.n512 VSS.n511 585
R252 VSS.n2108 VSS.n512 585
R253 VSS.n2106 VSS.n2105 585
R254 VSS.n2107 VSS.n2106 585
R255 VSS.n2104 VSS.n517 585
R256 VSS.n517 VSS.n516 585
R257 VSS.n788 VSS.n787 585
R258 VSS.n2013 VSS.n2012 585
R259 VSS.n2011 VSS.n799 585
R260 VSS.n2015 VSS.n799 585
R261 VSS.n2010 VSS.n2009 585
R262 VSS.n2008 VSS.n2007 585
R263 VSS.n2006 VSS.n2005 585
R264 VSS.n2004 VSS.n2003 585
R265 VSS.n2002 VSS.n2001 585
R266 VSS.n2000 VSS.n1999 585
R267 VSS.n1998 VSS.n1997 585
R268 VSS.n1996 VSS.n1995 585
R269 VSS.n1994 VSS.n1993 585
R270 VSS.n1992 VSS.n1991 585
R271 VSS.n1990 VSS.n1989 585
R272 VSS.n1988 VSS.n1987 585
R273 VSS.n1986 VSS.n1985 585
R274 VSS.n1984 VSS.n1983 585
R275 VSS.n1982 VSS.n1981 585
R276 VSS.n1980 VSS.n1979 585
R277 VSS.n1978 VSS.n798 585
R278 VSS.n2015 VSS.n798 585
R279 VSS.n1229 VSS.n1228 585
R280 VSS.n1227 VSS.n1226 585
R281 VSS.n1225 VSS.n1224 585
R282 VSS.n1223 VSS.n1222 585
R283 VSS.n1221 VSS.n1220 585
R284 VSS.n1219 VSS.n1218 585
R285 VSS.n1217 VSS.n1216 585
R286 VSS.n1215 VSS.n1214 585
R287 VSS.n1213 VSS.n1212 585
R288 VSS.n1211 VSS.n1210 585
R289 VSS.n1209 VSS.n1208 585
R290 VSS.n1207 VSS.n1206 585
R291 VSS.n1205 VSS.n1204 585
R292 VSS.n1203 VSS.n1202 585
R293 VSS.n1201 VSS.n1200 585
R294 VSS.n1199 VSS.n1198 585
R295 VSS.n1197 VSS.n1196 585
R296 VSS.n1195 VSS.n1194 585
R297 VSS.n1193 VSS.n1192 585
R298 VSS.n649 VSS.n647 585
R299 VSS.n2092 VSS.n2091 585
R300 VSS.n2093 VSS.n2092 585
R301 VSS.n2090 VSS.n648 585
R302 VSS.n648 VSS.n646 585
R303 VSS.n2089 VSS.n2088 585
R304 VSS.n2088 VSS.n2087 585
R305 VSS.n651 VSS.n650 585
R306 VSS.n2086 VSS.n651 585
R307 VSS.n2084 VSS.n2083 585
R308 VSS.n2085 VSS.n2084 585
R309 VSS.n2082 VSS.n653 585
R310 VSS.n653 VSS.n652 585
R311 VSS.n2081 VSS.n2080 585
R312 VSS.n2080 VSS.n2079 585
R313 VSS.n655 VSS.n654 585
R314 VSS.n2078 VSS.n655 585
R315 VSS.n2076 VSS.n2075 585
R316 VSS.n2077 VSS.n2076 585
R317 VSS.n2074 VSS.n657 585
R318 VSS.n657 VSS.n656 585
R319 VSS.n2073 VSS.n2072 585
R320 VSS.n2072 VSS.n2071 585
R321 VSS.n659 VSS.n658 585
R322 VSS.n2070 VSS.n659 585
R323 VSS.n2068 VSS.n2067 585
R324 VSS.n2069 VSS.n2068 585
R325 VSS.n2066 VSS.n661 585
R326 VSS.n661 VSS.n660 585
R327 VSS.n2065 VSS.n2064 585
R328 VSS.n2064 VSS.n2063 585
R329 VSS.n663 VSS.n662 585
R330 VSS.n2062 VSS.n663 585
R331 VSS.n2060 VSS.n2059 585
R332 VSS.n2061 VSS.n2060 585
R333 VSS.n2058 VSS.n665 585
R334 VSS.n1035 VSS.n665 585
R335 VSS.n1042 VSS.n667 585
R336 VSS.n1043 VSS.n1042 585
R337 VSS.n1041 VSS.n1040 585
R338 VSS.n1041 VSS.n1036 585
R339 VSS.n1039 VSS.n1038 585
R340 VSS.n1038 VSS.n1037 585
R341 VSS.n770 VSS.n769 585
R342 VSS.n772 VSS.n770 585
R343 VSS.n2050 VSS.n2049 585
R344 VSS.n2049 VSS.n2048 585
R345 VSS.n774 VSS.n771 585
R346 VSS.n2047 VSS.n771 585
R347 VSS.n2045 VSS.n2044 585
R348 VSS.n2046 VSS.n2045 585
R349 VSS.n2043 VSS.n773 585
R350 VSS.n777 VSS.n773 585
R351 VSS.n2042 VSS.n2041 585
R352 VSS.n2041 VSS.n2040 585
R353 VSS.n776 VSS.n775 585
R354 VSS.n2039 VSS.n776 585
R355 VSS.n2037 VSS.n2036 585
R356 VSS.n2038 VSS.n2037 585
R357 VSS.n2035 VSS.n778 585
R358 VSS.n781 VSS.n778 585
R359 VSS.n2034 VSS.n2033 585
R360 VSS.n2033 VSS.n2032 585
R361 VSS.n780 VSS.n779 585
R362 VSS.n2031 VSS.n780 585
R363 VSS.n2029 VSS.n2028 585
R364 VSS.n2030 VSS.n2029 585
R365 VSS.n2027 VSS.n782 585
R366 VSS.n785 VSS.n782 585
R367 VSS.n2026 VSS.n2025 585
R368 VSS.n2025 VSS.n2024 585
R369 VSS.n784 VSS.n783 585
R370 VSS.n2023 VSS.n784 585
R371 VSS.n2021 VSS.n2020 585
R372 VSS.n2022 VSS.n2021 585
R373 VSS.n2019 VSS.n786 585
R374 VSS.n789 VSS.n786 585
R375 VSS.n2018 VSS.n2017 585
R376 VSS.n2017 VSS.n2016 585
R377 VSS.n1538 VSS.n1537 585
R378 VSS.n1536 VSS.n1118 585
R379 VSS.n1535 VSS.n1117 585
R380 VSS.n1540 VSS.n1117 585
R381 VSS.n1534 VSS.n1533 585
R382 VSS.n1532 VSS.n1531 585
R383 VSS.n1530 VSS.n1529 585
R384 VSS.n1528 VSS.n1527 585
R385 VSS.n1526 VSS.n1525 585
R386 VSS.n1524 VSS.n1523 585
R387 VSS.n1522 VSS.n1521 585
R388 VSS.n1520 VSS.n1519 585
R389 VSS.n1518 VSS.n1517 585
R390 VSS.n1516 VSS.n1515 585
R391 VSS.n1514 VSS.n1513 585
R392 VSS.n1512 VSS.n1511 585
R393 VSS.n1510 VSS.n1509 585
R394 VSS.n1508 VSS.n1507 585
R395 VSS.n1506 VSS.n1505 585
R396 VSS.n1504 VSS.n1503 585
R397 VSS.n1502 VSS.n1501 585
R398 VSS.n1500 VSS.n1499 585
R399 VSS.n1498 VSS.n1497 585
R400 VSS.n1496 VSS.n1495 585
R401 VSS.n1494 VSS.n1121 585
R402 VSS.n1494 VSS.n1493 585
R403 VSS.n1471 VSS.n1122 585
R404 VSS.n1123 VSS.n1122 585
R405 VSS.n1472 VSS.n1131 585
R406 VSS.n1484 VSS.n1131 585
R407 VSS.n1474 VSS.n1139 585
R408 VSS.n1139 VSS.n1130 585
R409 VSS.n1476 VSS.n1475 585
R410 VSS.n1477 VSS.n1476 585
R411 VSS.n1469 VSS.n1138 585
R412 VSS.n1381 VSS.n1138 585
R413 VSS.n1468 VSS.n1467 585
R414 VSS.n1467 VSS.n1466 585
R415 VSS.n1141 VSS.n1140 585
R416 VSS.n1385 VSS.n1141 585
R417 VSS.n1459 VSS.n1458 585
R418 VSS.n1460 VSS.n1459 585
R419 VSS.n1457 VSS.n1147 585
R420 VSS.n1151 VSS.n1147 585
R421 VSS.n1456 VSS.n1455 585
R422 VSS.n1455 VSS.n1454 585
R423 VSS.n1149 VSS.n1148 585
R424 VSS.n1150 VSS.n1149 585
R425 VSS.n1411 VSS.n1410 585
R426 VSS.n1413 VSS.n1408 585
R427 VSS.n1415 VSS.n1414 585
R428 VSS.n1416 VSS.n1407 585
R429 VSS.n1418 VSS.n1417 585
R430 VSS.n1420 VSS.n1405 585
R431 VSS.n1422 VSS.n1421 585
R432 VSS.n1423 VSS.n1404 585
R433 VSS.n1425 VSS.n1424 585
R434 VSS.n1427 VSS.n1402 585
R435 VSS.n1429 VSS.n1428 585
R436 VSS.n1430 VSS.n1401 585
R437 VSS.n1432 VSS.n1431 585
R438 VSS.n1434 VSS.n1399 585
R439 VSS.n1436 VSS.n1435 585
R440 VSS.n1437 VSS.n1398 585
R441 VSS.n1439 VSS.n1438 585
R442 VSS.n1441 VSS.n1396 585
R443 VSS.n1443 VSS.n1442 585
R444 VSS.n1444 VSS.n1395 585
R445 VSS.n1446 VSS.n1445 585
R446 VSS.n1448 VSS.n1394 585
R447 VSS.n1450 VSS.n1449 585
R448 VSS.n1449 VSS.n98 585
R449 VSS.n1451 VSS.n1393 585
R450 VSS.n1393 VSS.n1150 585
R451 VSS.n1453 VSS.n1452 585
R452 VSS.n1454 VSS.n1453 585
R453 VSS.n1145 VSS.n1144 585
R454 VSS.n1151 VSS.n1145 585
R455 VSS.n1462 VSS.n1461 585
R456 VSS.n1461 VSS.n1460 585
R457 VSS.n1463 VSS.n1143 585
R458 VSS.n1385 VSS.n1143 585
R459 VSS.n1465 VSS.n1464 585
R460 VSS.n1466 VSS.n1465 585
R461 VSS.n1136 VSS.n1135 585
R462 VSS.n1381 VSS.n1136 585
R463 VSS.n1479 VSS.n1478 585
R464 VSS.n1478 VSS.n1477 585
R465 VSS.n1480 VSS.n1133 585
R466 VSS.n1133 VSS.n1130 585
R467 VSS.n1483 VSS.n1482 585
R468 VSS.n1484 VSS.n1483 585
R469 VSS.n1481 VSS.n1134 585
R470 VSS.n1134 VSS.n1123 585
R471 VSS.n1120 VSS.n1119 585
R472 VSS.n1493 VSS.n1119 585
R473 VSS.n1815 VSS.n856 585
R474 VSS.n1814 VSS.n1813 585
R475 VSS.n1811 VSS.n858 585
R476 VSS.n1811 VSS.n855 585
R477 VSS.n1810 VSS.n1809 585
R478 VSS.n1808 VSS.n1807 585
R479 VSS.n1806 VSS.n860 585
R480 VSS.n1804 VSS.n1803 585
R481 VSS.n1802 VSS.n861 585
R482 VSS.n1801 VSS.n1800 585
R483 VSS.n1798 VSS.n862 585
R484 VSS.n1796 VSS.n1795 585
R485 VSS.n1792 VSS.n863 585
R486 VSS.n1791 VSS.n1790 585
R487 VSS.n1788 VSS.n865 585
R488 VSS.n1786 VSS.n1785 585
R489 VSS.n1784 VSS.n866 585
R490 VSS.n1783 VSS.n1782 585
R491 VSS.n1780 VSS.n867 585
R492 VSS.n1778 VSS.n1777 585
R493 VSS.n1776 VSS.n868 585
R494 VSS.n1775 VSS.n1774 585
R495 VSS.n1772 VSS.n869 585
R496 VSS.n1770 VSS.n1769 585
R497 VSS.n1768 VSS.n854 585
R498 VSS.n1818 VSS.n854 585
R499 VSS.n1767 VSS.n853 585
R500 VSS.n1819 VSS.n853 585
R501 VSS.n1766 VSS.n852 585
R502 VSS.n1820 VSS.n852 585
R503 VSS.n1765 VSS.n1764 585
R504 VSS.n1764 VSS.n840 585
R505 VSS.n1763 VSS.n839 585
R506 VSS.n1974 VSS.n839 585
R507 VSS.n1762 VSS.n1761 585
R508 VSS.n1761 VSS.n802 585
R509 VSS.n1760 VSS.n846 585
R510 VSS.n1828 VSS.n846 585
R511 VSS.n1759 VSS.n1758 585
R512 VSS.n1758 VSS.n1757 585
R513 VSS.n1756 VSS.n870 585
R514 VSS.n1756 VSS.n1755 585
R515 VSS.n1687 VSS.n871 585
R516 VSS.n879 VSS.n871 585
R517 VSS.n1688 VSS.n878 585
R518 VSS.n1749 VSS.n878 585
R519 VSS.n1691 VSS.n1689 585
R520 VSS.n1691 VSS.n1690 585
R521 VSS.n1693 VSS.n1692 585
R522 VSS.n1695 VSS.n1694 585
R523 VSS.n1697 VSS.n1696 585
R524 VSS.n1699 VSS.n1698 585
R525 VSS.n1701 VSS.n1700 585
R526 VSS.n1703 VSS.n1702 585
R527 VSS.n1705 VSS.n1704 585
R528 VSS.n1707 VSS.n1706 585
R529 VSS.n1709 VSS.n1708 585
R530 VSS.n1711 VSS.n1710 585
R531 VSS.n1713 VSS.n1712 585
R532 VSS.n1715 VSS.n1714 585
R533 VSS.n1717 VSS.n1716 585
R534 VSS.n1719 VSS.n1718 585
R535 VSS.n1721 VSS.n1720 585
R536 VSS.n1723 VSS.n1722 585
R537 VSS.n1725 VSS.n1724 585
R538 VSS.n1727 VSS.n1726 585
R539 VSS.n1729 VSS.n1728 585
R540 VSS.n1731 VSS.n1730 585
R541 VSS.n1733 VSS.n1732 585
R542 VSS.n1734 VSS.n1686 585
R543 VSS.n1736 VSS.n1735 585
R544 VSS.n1737 VSS.n1736 585
R545 VSS.n876 VSS.n875 585
R546 VSS.n1690 VSS.n876 585
R547 VSS.n1751 VSS.n1750 585
R548 VSS.n1750 VSS.n1749 585
R549 VSS.n1752 VSS.n874 585
R550 VSS.n879 VSS.n874 585
R551 VSS.n1754 VSS.n1753 585
R552 VSS.n1755 VSS.n1754 585
R553 VSS.n849 VSS.n847 585
R554 VSS.n1757 VSS.n847 585
R555 VSS.n1827 VSS.n1826 585
R556 VSS.n1828 VSS.n1827 585
R557 VSS.n1825 VSS.n848 585
R558 VSS.n848 VSS.n802 585
R559 VSS.n1824 VSS.n841 585
R560 VSS.n1974 VSS.n841 585
R561 VSS.n1823 VSS.n1822 585
R562 VSS.n1822 VSS.n840 585
R563 VSS.n1821 VSS.n850 585
R564 VSS.n1821 VSS.n1820 585
R565 VSS.n857 VSS.n851 585
R566 VSS.n1819 VSS.n851 585
R567 VSS.n1817 VSS.n1816 585
R568 VSS.n1818 VSS.n1817 585
R569 VSS.n2448 VSS.n2447 585
R570 VSS.n2446 VSS.n100 585
R571 VSS.n2445 VSS.n99 585
R572 VSS.n2450 VSS.n99 585
R573 VSS.n2444 VSS.n2443 585
R574 VSS.n2442 VSS.n2441 585
R575 VSS.n2440 VSS.n2439 585
R576 VSS.n2438 VSS.n2437 585
R577 VSS.n2436 VSS.n2435 585
R578 VSS.n2434 VSS.n2433 585
R579 VSS.n2432 VSS.n2431 585
R580 VSS.n2430 VSS.n2429 585
R581 VSS.n2428 VSS.n2427 585
R582 VSS.n2426 VSS.n2425 585
R583 VSS.n2424 VSS.n2423 585
R584 VSS.n2422 VSS.n2421 585
R585 VSS.n2420 VSS.n2419 585
R586 VSS.n2418 VSS.n2417 585
R587 VSS.n2416 VSS.n2415 585
R588 VSS.n2414 VSS.n2413 585
R589 VSS.n2412 VSS.n2411 585
R590 VSS.n2402 VSS.n2401 585
R591 VSS.n2404 VSS.n2403 585
R592 VSS.n2407 VSS.n2406 585
R593 VSS.n79 VSS.n76 585
R594 VSS.n2453 VSS.n2452 585
R595 VSS.n78 VSS.n77 585
R596 VSS.n2369 VSS.n2368 585
R597 VSS.n2371 VSS.n2370 585
R598 VSS.n2373 VSS.n2372 585
R599 VSS.n2375 VSS.n2374 585
R600 VSS.n2377 VSS.n2376 585
R601 VSS.n2379 VSS.n2378 585
R602 VSS.n2381 VSS.n2380 585
R603 VSS.n2383 VSS.n2382 585
R604 VSS.n2385 VSS.n2384 585
R605 VSS.n2387 VSS.n2386 585
R606 VSS.n2389 VSS.n2388 585
R607 VSS.n2391 VSS.n2390 585
R608 VSS.n2393 VSS.n2392 585
R609 VSS.n2394 VSS.n106 585
R610 VSS.n106 VSS.n80 585
R611 VSS.n2396 VSS.n2395 585
R612 VSS.n2397 VSS.n2396 585
R613 VSS.n2367 VSS.n105 585
R614 VSS.n105 VSS.n104 585
R615 VSS.n2366 VSS.n2365 585
R616 VSS.n2365 VSS.n2364 585
R617 VSS.n108 VSS.n107 585
R618 VSS.n109 VSS.n108 585
R619 VSS.n2357 VSS.n2356 585
R620 VSS.n2358 VSS.n2357 585
R621 VSS.n2355 VSS.n113 585
R622 VSS.n117 VSS.n113 585
R623 VSS.n2354 VSS.n2353 585
R624 VSS.n2353 VSS.n2352 585
R625 VSS.n115 VSS.n114 585
R626 VSS.n116 VSS.n115 585
R627 VSS.n2345 VSS.n2344 585
R628 VSS.n2346 VSS.n2345 585
R629 VSS.n2343 VSS.n121 585
R630 VSS.n125 VSS.n121 585
R631 VSS.n2342 VSS.n2341 585
R632 VSS.n2341 VSS.n2340 585
R633 VSS.n123 VSS.n122 585
R634 VSS.n124 VSS.n123 585
R635 VSS.n2333 VSS.n2332 585
R636 VSS.n2334 VSS.n2333 585
R637 VSS.n2331 VSS.n129 585
R638 VSS.n133 VSS.n129 585
R639 VSS.n2330 VSS.n2329 585
R640 VSS.n2329 VSS.n2328 585
R641 VSS.n131 VSS.n130 585
R642 VSS.n132 VSS.n131 585
R643 VSS.n2321 VSS.n2320 585
R644 VSS.n2322 VSS.n2321 585
R645 VSS.n2319 VSS.n137 585
R646 VSS.n141 VSS.n137 585
R647 VSS.n2318 VSS.n2317 585
R648 VSS.n2317 VSS.n2316 585
R649 VSS.n139 VSS.n138 585
R650 VSS.n140 VSS.n139 585
R651 VSS.n2309 VSS.n2308 585
R652 VSS.n2310 VSS.n2309 585
R653 VSS.n2307 VSS.n145 585
R654 VSS.n149 VSS.n145 585
R655 VSS.n2306 VSS.n2305 585
R656 VSS.n2305 VSS.n2304 585
R657 VSS.n147 VSS.n146 585
R658 VSS.n148 VSS.n147 585
R659 VSS.n2297 VSS.n2296 585
R660 VSS.n2298 VSS.n2297 585
R661 VSS.n2295 VSS.n154 585
R662 VSS.n154 VSS.n153 585
R663 VSS.n2294 VSS.n2293 585
R664 VSS.n2293 VSS.n2292 585
R665 VSS.n156 VSS.n155 585
R666 VSS.n157 VSS.n156 585
R667 VSS.n2285 VSS.n2284 585
R668 VSS.n2286 VSS.n2285 585
R669 VSS.n2283 VSS.n162 585
R670 VSS.n162 VSS.n161 585
R671 VSS.n2282 VSS.n2281 585
R672 VSS.n2281 VSS.n2280 585
R673 VSS.n164 VSS.n163 585
R674 VSS.n165 VSS.n164 585
R675 VSS.n2273 VSS.n2272 585
R676 VSS.n2274 VSS.n2273 585
R677 VSS.n2271 VSS.n170 585
R678 VSS.n170 VSS.n169 585
R679 VSS.n2270 VSS.n2269 585
R680 VSS.n2269 VSS.n2268 585
R681 VSS.n172 VSS.n171 585
R682 VSS.n173 VSS.n172 585
R683 VSS.n2261 VSS.n2260 585
R684 VSS.n2262 VSS.n2261 585
R685 VSS.n2259 VSS.n178 585
R686 VSS.n178 VSS.n177 585
R687 VSS.n2258 VSS.n2257 585
R688 VSS.n2257 VSS.n2256 585
R689 VSS.n180 VSS.n179 585
R690 VSS.n2249 VSS.n180 585
R691 VSS.n2248 VSS.n2247 585
R692 VSS.n2250 VSS.n2248 585
R693 VSS.n2246 VSS.n185 585
R694 VSS.n185 VSS.n184 585
R695 VSS.n2245 VSS.n2244 585
R696 VSS.n2244 VSS.n2243 585
R697 VSS.n187 VSS.n186 585
R698 VSS.n2236 VSS.n187 585
R699 VSS.n2235 VSS.n2234 585
R700 VSS.n2237 VSS.n2235 585
R701 VSS.n2233 VSS.n192 585
R702 VSS.n192 VSS.n191 585
R703 VSS.n2232 VSS.n2231 585
R704 VSS.n2231 VSS.n2230 585
R705 VSS.n194 VSS.n193 585
R706 VSS.n2223 VSS.n194 585
R707 VSS.n2222 VSS.n2221 585
R708 VSS.n2224 VSS.n2222 585
R709 VSS.n2220 VSS.n199 585
R710 VSS.n199 VSS.n198 585
R711 VSS.n2219 VSS.n2218 585
R712 VSS.n2218 VSS.n2217 585
R713 VSS.n201 VSS.n200 585
R714 VSS.n2210 VSS.n201 585
R715 VSS.n2209 VSS.n2208 585
R716 VSS.n2211 VSS.n2209 585
R717 VSS.n2207 VSS.n206 585
R718 VSS.n206 VSS.n205 585
R719 VSS.n2206 VSS.n2205 585
R720 VSS.n2205 VSS.n2204 585
R721 VSS.n208 VSS.n207 585
R722 VSS.n2196 VSS.n208 585
R723 VSS.n434 VSS.n433 585
R724 VSS.n2198 VSS.n434 585
R725 VSS.n432 VSS.n213 585
R726 VSS.n213 VSS.n212 585
R727 VSS.n431 VSS.n430 585
R728 VSS.n430 VSS.n429 585
R729 VSS.n215 VSS.n214 585
R730 VSS.n216 VSS.n215 585
R731 VSS.n422 VSS.n421 585
R732 VSS.n423 VSS.n422 585
R733 VSS.n420 VSS.n221 585
R734 VSS.n419 VSS.n418 585
R735 VSS.n416 VSS.n222 585
R736 VSS.n414 VSS.n413 585
R737 VSS.n412 VSS.n223 585
R738 VSS.n411 VSS.n410 585
R739 VSS.n408 VSS.n224 585
R740 VSS.n406 VSS.n405 585
R741 VSS.n404 VSS.n225 585
R742 VSS.n403 VSS.n402 585
R743 VSS.n400 VSS.n226 585
R744 VSS.n398 VSS.n397 585
R745 VSS.n396 VSS.n227 585
R746 VSS.n395 VSS.n394 585
R747 VSS.n392 VSS.n228 585
R748 VSS.n390 VSS.n389 585
R749 VSS.n230 VSS.n229 585
R750 VSS.n284 VSS.n283 585
R751 VSS.n281 VSS.n232 585
R752 VSS.n279 VSS.n278 585
R753 VSS.n277 VSS.n233 585
R754 VSS.n276 VSS.n275 585
R755 VSS.n273 VSS.n234 585
R756 VSS.n271 VSS.n270 585
R757 VSS.n269 VSS.n235 585
R758 VSS.n268 VSS.n267 585
R759 VSS.n265 VSS.n236 585
R760 VSS.n263 VSS.n262 585
R761 VSS.n261 VSS.n237 585
R762 VSS.n260 VSS.n259 585
R763 VSS.n257 VSS.n238 585
R764 VSS.n255 VSS.n254 585
R765 VSS.n253 VSS.n239 585
R766 VSS.n252 VSS.n251 585
R767 VSS.n249 VSS.n240 585
R768 VSS.n247 VSS.n246 585
R769 VSS.n245 VSS.n241 585
R770 VSS.n244 VSS.n243 585
R771 VSS.n219 VSS.n218 585
R772 VSS.n220 VSS.n219 585
R773 VSS.n425 VSS.n424 585
R774 VSS.n424 VSS.n423 585
R775 VSS.n426 VSS.n217 585
R776 VSS.n217 VSS.n216 585
R777 VSS.n428 VSS.n427 585
R778 VSS.n429 VSS.n428 585
R779 VSS.n211 VSS.n210 585
R780 VSS.n212 VSS.n211 585
R781 VSS.n2200 VSS.n2199 585
R782 VSS.n2199 VSS.n2198 585
R783 VSS.n2201 VSS.n209 585
R784 VSS.n2196 VSS.n209 585
R785 VSS.n2203 VSS.n2202 585
R786 VSS.n2204 VSS.n2203 585
R787 VSS.n204 VSS.n203 585
R788 VSS.n205 VSS.n204 585
R789 VSS.n2213 VSS.n2212 585
R790 VSS.n2212 VSS.n2211 585
R791 VSS.n2214 VSS.n202 585
R792 VSS.n2210 VSS.n202 585
R793 VSS.n2216 VSS.n2215 585
R794 VSS.n2217 VSS.n2216 585
R795 VSS.n197 VSS.n196 585
R796 VSS.n198 VSS.n197 585
R797 VSS.n2226 VSS.n2225 585
R798 VSS.n2225 VSS.n2224 585
R799 VSS.n2227 VSS.n195 585
R800 VSS.n2223 VSS.n195 585
R801 VSS.n2229 VSS.n2228 585
R802 VSS.n2230 VSS.n2229 585
R803 VSS.n190 VSS.n189 585
R804 VSS.n191 VSS.n190 585
R805 VSS.n2239 VSS.n2238 585
R806 VSS.n2238 VSS.n2237 585
R807 VSS.n2240 VSS.n188 585
R808 VSS.n2236 VSS.n188 585
R809 VSS.n2242 VSS.n2241 585
R810 VSS.n2243 VSS.n2242 585
R811 VSS.n183 VSS.n182 585
R812 VSS.n184 VSS.n183 585
R813 VSS.n2252 VSS.n2251 585
R814 VSS.n2251 VSS.n2250 585
R815 VSS.n2253 VSS.n181 585
R816 VSS.n2249 VSS.n181 585
R817 VSS.n2255 VSS.n2254 585
R818 VSS.n2256 VSS.n2255 585
R819 VSS.n176 VSS.n175 585
R820 VSS.n177 VSS.n176 585
R821 VSS.n2264 VSS.n2263 585
R822 VSS.n2263 VSS.n2262 585
R823 VSS.n2265 VSS.n174 585
R824 VSS.n174 VSS.n173 585
R825 VSS.n2267 VSS.n2266 585
R826 VSS.n2268 VSS.n2267 585
R827 VSS.n168 VSS.n167 585
R828 VSS.n169 VSS.n168 585
R829 VSS.n2276 VSS.n2275 585
R830 VSS.n2275 VSS.n2274 585
R831 VSS.n2277 VSS.n166 585
R832 VSS.n166 VSS.n165 585
R833 VSS.n2279 VSS.n2278 585
R834 VSS.n2280 VSS.n2279 585
R835 VSS.n160 VSS.n159 585
R836 VSS.n161 VSS.n160 585
R837 VSS.n2288 VSS.n2287 585
R838 VSS.n2287 VSS.n2286 585
R839 VSS.n2289 VSS.n158 585
R840 VSS.n158 VSS.n157 585
R841 VSS.n2291 VSS.n2290 585
R842 VSS.n2292 VSS.n2291 585
R843 VSS.n152 VSS.n151 585
R844 VSS.n153 VSS.n152 585
R845 VSS.n2300 VSS.n2299 585
R846 VSS.n2299 VSS.n2298 585
R847 VSS.n2301 VSS.n150 585
R848 VSS.n150 VSS.n148 585
R849 VSS.n2303 VSS.n2302 585
R850 VSS.n2304 VSS.n2303 585
R851 VSS.n144 VSS.n143 585
R852 VSS.n149 VSS.n144 585
R853 VSS.n2312 VSS.n2311 585
R854 VSS.n2311 VSS.n2310 585
R855 VSS.n2313 VSS.n142 585
R856 VSS.n142 VSS.n140 585
R857 VSS.n2315 VSS.n2314 585
R858 VSS.n2316 VSS.n2315 585
R859 VSS.n136 VSS.n135 585
R860 VSS.n141 VSS.n136 585
R861 VSS.n2324 VSS.n2323 585
R862 VSS.n2323 VSS.n2322 585
R863 VSS.n2325 VSS.n134 585
R864 VSS.n134 VSS.n132 585
R865 VSS.n2327 VSS.n2326 585
R866 VSS.n2328 VSS.n2327 585
R867 VSS.n128 VSS.n127 585
R868 VSS.n133 VSS.n128 585
R869 VSS.n2336 VSS.n2335 585
R870 VSS.n2335 VSS.n2334 585
R871 VSS.n2337 VSS.n126 585
R872 VSS.n126 VSS.n124 585
R873 VSS.n2339 VSS.n2338 585
R874 VSS.n2340 VSS.n2339 585
R875 VSS.n120 VSS.n119 585
R876 VSS.n125 VSS.n120 585
R877 VSS.n2348 VSS.n2347 585
R878 VSS.n2347 VSS.n2346 585
R879 VSS.n2349 VSS.n118 585
R880 VSS.n118 VSS.n116 585
R881 VSS.n2351 VSS.n2350 585
R882 VSS.n2352 VSS.n2351 585
R883 VSS.n112 VSS.n111 585
R884 VSS.n117 VSS.n112 585
R885 VSS.n2360 VSS.n2359 585
R886 VSS.n2359 VSS.n2358 585
R887 VSS.n2361 VSS.n110 585
R888 VSS.n110 VSS.n109 585
R889 VSS.n2363 VSS.n2362 585
R890 VSS.n2364 VSS.n2363 585
R891 VSS.n103 VSS.n102 585
R892 VSS.n104 VSS.n103 585
R893 VSS.n2399 VSS.n2398 585
R894 VSS.n2398 VSS.n2397 585
R895 VSS.n2400 VSS.n101 585
R896 VSS.n101 VSS.n80 585
R897 VSS.n1977 VSS.n1976 585
R898 VSS.n801 VSS.n800 585
R899 VSS.n1973 VSS.n1972 585
R900 VSS.n1974 VSS.n1973 585
R901 VSS.n1971 VSS.n842 585
R902 VSS.n1970 VSS.n1969 585
R903 VSS.n1968 VSS.n1967 585
R904 VSS.n1966 VSS.n1965 585
R905 VSS.n1964 VSS.n1963 585
R906 VSS.n1962 VSS.n1961 585
R907 VSS.n1960 VSS.n1959 585
R908 VSS.n1958 VSS.n1957 585
R909 VSS.n1956 VSS.n1955 585
R910 VSS.n1954 VSS.n1953 585
R911 VSS.n1952 VSS.n1951 585
R912 VSS.n1950 VSS.n1949 585
R913 VSS.n1948 VSS.n1947 585
R914 VSS.n1946 VSS.n1945 585
R915 VSS.n1944 VSS.n1943 585
R916 VSS.n1942 VSS.n1941 585
R917 VSS.n1940 VSS.n1939 585
R918 VSS.n1938 VSS.n1937 585
R919 VSS.n1936 VSS.n1935 585
R920 VSS.n1934 VSS.n1933 585
R921 VSS.n1932 VSS.n1931 585
R922 VSS.n1930 VSS.n1929 585
R923 VSS.n1928 VSS.n1927 585
R924 VSS.n1926 VSS.n1925 585
R925 VSS.n1924 VSS.n1923 585
R926 VSS.n1922 VSS.n1921 585
R927 VSS.n1920 VSS.n1919 585
R928 VSS.n1918 VSS.n1917 585
R929 VSS.n1916 VSS.n1915 585
R930 VSS.n1914 VSS.n1913 585
R931 VSS.n1912 VSS.n1911 585
R932 VSS.n1910 VSS.n1909 585
R933 VSS.n1908 VSS.n1907 585
R934 VSS.n1906 VSS.n1905 585
R935 VSS.n1904 VSS.n1903 585
R936 VSS.n1902 VSS.n1901 585
R937 VSS.n1900 VSS.n1899 585
R938 VSS.n1898 VSS.n1897 585
R939 VSS.n1896 VSS.n1895 585
R940 VSS.n1894 VSS.n1893 585
R941 VSS.n1892 VSS.n1891 585
R942 VSS.n1890 VSS.n1889 585
R943 VSS.n1888 VSS.n1887 585
R944 VSS.n1886 VSS.n1885 585
R945 VSS.n1884 VSS.n1883 585
R946 VSS.n1882 VSS.n1881 585
R947 VSS.n1880 VSS.n1879 585
R948 VSS.n1878 VSS.n1877 585
R949 VSS.n1876 VSS.n1875 585
R950 VSS.n1874 VSS.n1873 585
R951 VSS.n1872 VSS.n1871 585
R952 VSS.n1870 VSS.n1869 585
R953 VSS.n1868 VSS.n1867 585
R954 VSS.n1866 VSS.n1865 585
R955 VSS.n1864 VSS.n1863 585
R956 VSS.n1862 VSS.n1861 585
R957 VSS.n1860 VSS.n1859 585
R958 VSS.n1858 VSS.n1857 585
R959 VSS.n1856 VSS.n1855 585
R960 VSS.n1854 VSS.n1853 585
R961 VSS.n1852 VSS.n1851 585
R962 VSS.n1850 VSS.n1849 585
R963 VSS.n1848 VSS.n1847 585
R964 VSS.n1846 VSS.n1845 585
R965 VSS.n1844 VSS.n1843 585
R966 VSS.n1842 VSS.n1841 585
R967 VSS.n1840 VSS.n1839 585
R968 VSS.n1838 VSS.n1837 585
R969 VSS.n1836 VSS.n1835 585
R970 VSS.n1834 VSS.n1833 585
R971 VSS.n1832 VSS.n838 585
R972 VSS.n1974 VSS.n838 585
R973 VSS.n1831 VSS.n1830 585
R974 VSS.n1830 VSS.n1829 585
R975 VSS.n844 VSS.n843 585
R976 VSS.n845 VSS.n844 585
R977 VSS.n1744 VSS.n1743 585
R978 VSS.n1743 VSS.n873 585
R979 VSS.n1745 VSS.n881 585
R980 VSS.n881 VSS.n872 585
R981 VSS.n1747 VSS.n1746 585
R982 VSS.n1748 VSS.n1747 585
R983 VSS.n1742 VSS.n880 585
R984 VSS.n880 VSS.n877 585
R985 VSS.n1741 VSS.n1740 585
R986 VSS.n1740 VSS.n1739 585
R987 VSS.n883 VSS.n882 585
R988 VSS.n1738 VSS.n883 585
R989 VSS.n1673 VSS.n1672 585
R990 VSS.n1674 VSS.n1673 585
R991 VSS.n1671 VSS.n885 585
R992 VSS.n885 VSS.n884 585
R993 VSS.n1670 VSS.n1669 585
R994 VSS.n1669 VSS.n1668 585
R995 VSS.n887 VSS.n886 585
R996 VSS.n888 VSS.n887 585
R997 VSS.n1618 VSS.n1617 585
R998 VSS.n1619 VSS.n1618 585
R999 VSS.n1616 VSS.n907 585
R1000 VSS.n907 VSS.n906 585
R1001 VSS.n1615 VSS.n1614 585
R1002 VSS.n1614 VSS.n1613 585
R1003 VSS.n909 VSS.n908 585
R1004 VSS.n1604 VSS.n909 585
R1005 VSS.n1578 VSS.n1577 585
R1006 VSS.n1578 VSS.n916 585
R1007 VSS.n1582 VSS.n1581 585
R1008 VSS.n1581 VSS.n1580 585
R1009 VSS.n1583 VSS.n929 585
R1010 VSS.n929 VSS.n921 585
R1011 VSS.n1585 VSS.n1584 585
R1012 VSS.n1586 VSS.n1585 585
R1013 VSS.n930 VSS.n928 585
R1014 VSS.n928 VSS.n925 585
R1015 VSS.n1568 VSS.n1567 585
R1016 VSS.n1567 VSS.n1566 585
R1017 VSS.n1034 VSS.n1033 585
R1018 VSS.n1048 VSS.n1034 585
R1019 VSS.n1546 VSS.n1103 585
R1020 VSS.n1103 VSS.n1047 585
R1021 VSS.n1548 VSS.n1547 585
R1022 VSS.n1549 VSS.n1548 585
R1023 VSS.n1545 VSS.n1102 585
R1024 VSS.n1541 VSS.n1102 585
R1025 VSS.n1544 VSS.n1543 585
R1026 VSS.n1543 VSS.n1542 585
R1027 VSS.n1105 VSS.n1104 585
R1028 VSS.n1106 VSS.n1105 585
R1029 VSS.n1489 VSS.n1126 585
R1030 VSS.n1126 VSS.n1125 585
R1031 VSS.n1491 VSS.n1490 585
R1032 VSS.n1492 VSS.n1491 585
R1033 VSS.n1488 VSS.n1124 585
R1034 VSS.n1132 VSS.n1124 585
R1035 VSS.n1487 VSS.n1486 585
R1036 VSS.n1486 VSS.n1485 585
R1037 VSS.n1128 VSS.n1127 585
R1038 VSS.n1129 VSS.n1128 585
R1039 VSS.n1379 VSS.n1378 585
R1040 VSS.n1378 VSS.n1137 585
R1041 VSS.n1383 VSS.n1380 585
R1042 VSS.n1383 VSS.n1382 585
R1043 VSS.n1384 VSS.n1377 585
R1044 VSS.n1384 VSS.n1142 585
R1045 VSS.n1388 VSS.n1387 585
R1046 VSS.n1387 VSS.n1386 585
R1047 VSS.n1389 VSS.n1153 585
R1048 VSS.n1153 VSS.n1146 585
R1049 VSS.n1391 VSS.n1390 585
R1050 VSS.n1392 VSS.n1391 585
R1051 VSS.n1376 VSS.n1152 585
R1052 VSS.n1375 VSS.n1374 585
R1053 VSS.n1155 VSS.n1154 585
R1054 VSS.n1370 VSS.n1369 585
R1055 VSS.n1368 VSS.n1191 585
R1056 VSS.n1367 VSS.n1366 585
R1057 VSS.n1365 VSS.n1364 585
R1058 VSS.n1363 VSS.n1362 585
R1059 VSS.n1361 VSS.n1360 585
R1060 VSS.n1359 VSS.n1358 585
R1061 VSS.n1357 VSS.n1356 585
R1062 VSS.n1355 VSS.n1354 585
R1063 VSS.n1353 VSS.n1352 585
R1064 VSS.n1351 VSS.n1350 585
R1065 VSS.n1349 VSS.n1348 585
R1066 VSS.n1347 VSS.n1346 585
R1067 VSS.n1345 VSS.n1344 585
R1068 VSS.n1343 VSS.n1342 585
R1069 VSS.n1341 VSS.n1340 585
R1070 VSS.n1339 VSS.n1338 585
R1071 VSS.n1337 VSS.n1336 585
R1072 VSS.n1335 VSS.n1334 585
R1073 VSS.n1333 VSS.n1332 585
R1074 VSS.n1331 VSS.n1330 585
R1075 VSS.n1329 VSS.n1328 585
R1076 VSS.n1327 VSS.n1326 585
R1077 VSS.n1325 VSS.n1324 585
R1078 VSS.n1323 VSS.n1322 585
R1079 VSS.n1321 VSS.n1320 585
R1080 VSS.n1319 VSS.n1318 585
R1081 VSS.n1317 VSS.n1316 585
R1082 VSS.n1315 VSS.n1314 585
R1083 VSS.n1313 VSS.n1312 585
R1084 VSS.n1311 VSS.n1310 585
R1085 VSS.n1309 VSS.n1308 585
R1086 VSS.n1307 VSS.n1306 585
R1087 VSS.n1305 VSS.n1304 585
R1088 VSS.n1303 VSS.n1302 585
R1089 VSS.n1301 VSS.n1300 585
R1090 VSS.n1299 VSS.n1298 585
R1091 VSS.n1297 VSS.n1296 585
R1092 VSS.n1295 VSS.n1294 585
R1093 VSS.n1293 VSS.n1292 585
R1094 VSS.n1291 VSS.n1290 585
R1095 VSS.n1289 VSS.n1288 585
R1096 VSS.n1287 VSS.n1286 585
R1097 VSS.n1285 VSS.n1284 585
R1098 VSS.n1283 VSS.n1282 585
R1099 VSS.n1281 VSS.n1280 585
R1100 VSS.n1279 VSS.n1278 585
R1101 VSS.n1277 VSS.n1276 585
R1102 VSS.n1275 VSS.n1274 585
R1103 VSS.n1273 VSS.n1272 585
R1104 VSS.n1271 VSS.n1270 585
R1105 VSS.n1269 VSS.n1268 585
R1106 VSS.n1267 VSS.n1266 585
R1107 VSS.n1265 VSS.n1264 585
R1108 VSS.n1263 VSS.n1262 585
R1109 VSS.n1261 VSS.n1260 585
R1110 VSS.n1259 VSS.n1258 585
R1111 VSS.n1257 VSS.n1256 585
R1112 VSS.n1255 VSS.n1254 585
R1113 VSS.n1253 VSS.n1252 585
R1114 VSS.n1251 VSS.n1250 585
R1115 VSS.n1249 VSS.n1248 585
R1116 VSS.n1247 VSS.n1246 585
R1117 VSS.n1245 VSS.n1244 585
R1118 VSS.n1243 VSS.n1242 585
R1119 VSS.n1241 VSS.n1240 585
R1120 VSS.n1239 VSS.n1238 585
R1121 VSS.n1237 VSS.n1236 585
R1122 VSS.n1235 VSS.n1234 585
R1123 VSS.n1233 VSS.n1232 585
R1124 VSS.n1231 VSS.n1230 585
R1125 VSS.n1046 VSS.n1045 585
R1126 VSS.n1550 VSS.n1046 585
R1127 VSS.n1100 VSS.n1099 585
R1128 VSS.n1098 VSS.n1063 585
R1129 VSS.n1097 VSS.n1096 585
R1130 VSS.n1095 VSS.n1094 585
R1131 VSS.n1093 VSS.n1092 585
R1132 VSS.n1091 VSS.n1090 585
R1133 VSS.n1089 VSS.n1088 585
R1134 VSS.n1087 VSS.n1086 585
R1135 VSS.n1085 VSS.n1084 585
R1136 VSS.n1083 VSS.n1082 585
R1137 VSS.n1081 VSS.n1080 585
R1138 VSS.n1079 VSS.n1078 585
R1139 VSS.n1077 VSS.n1076 585
R1140 VSS.n1075 VSS.n1074 585
R1141 VSS.n1073 VSS.n1072 585
R1142 VSS.n1071 VSS.n1070 585
R1143 VSS.n1069 VSS.n1068 585
R1144 VSS.n1067 VSS.n1066 585
R1145 VSS.n1065 VSS.n1064 585
R1146 VSS.n1053 VSS.n1052 585
R1147 VSS.n1553 VSS.n1552 585
R1148 VSS.n1554 VSS.n1049 585
R1149 VSS.n1557 VSS.n1556 585
R1150 VSS.n1558 VSS.n1557 585
R1151 VSS.n1555 VSS.n1051 585
R1152 VSS.n1051 VSS.n1050 585
R1153 VSS.n924 VSS.n923 585
R1154 VSS.n1565 VSS.n924 585
R1155 VSS.n1589 VSS.n1588 585
R1156 VSS.n1588 VSS.n1587 585
R1157 VSS.n1590 VSS.n922 585
R1158 VSS.n927 VSS.n922 585
R1159 VSS.n1592 VSS.n1591 585
R1160 VSS.n1593 VSS.n1592 585
R1161 VSS.n915 VSS.n914 585
R1162 VSS.n1579 VSS.n915 585
R1163 VSS.n1607 VSS.n1606 585
R1164 VSS.n1606 VSS.n1605 585
R1165 VSS.n1608 VSS.n912 585
R1166 VSS.n912 VSS.n910 585
R1167 VSS.n1611 VSS.n1610 585
R1168 VSS.n1612 VSS.n1611 585
R1169 VSS.n1609 VSS.n913 585
R1170 VSS.n913 VSS.n905 585
R1171 VSS.n902 VSS.n901 585
R1172 VSS.n1620 VSS.n901 585
R1173 VSS.n1665 VSS.n1664 585
R1174 VSS.n1663 VSS.n900 585
R1175 VSS.n1662 VSS.n899 585
R1176 VSS.n1667 VSS.n899 585
R1177 VSS.n1661 VSS.n1660 585
R1178 VSS.n1659 VSS.n1658 585
R1179 VSS.n1657 VSS.n1656 585
R1180 VSS.n1655 VSS.n1654 585
R1181 VSS.n1653 VSS.n1652 585
R1182 VSS.n1651 VSS.n1650 585
R1183 VSS.n1649 VSS.n1648 585
R1184 VSS.n1647 VSS.n1646 585
R1185 VSS.n1645 VSS.n1644 585
R1186 VSS.n1643 VSS.n1642 585
R1187 VSS.n1641 VSS.n1640 585
R1188 VSS.n1639 VSS.n1638 585
R1189 VSS.n1637 VSS.n1636 585
R1190 VSS.n1635 VSS.n1634 585
R1191 VSS.n1633 VSS.n1632 585
R1192 VSS.n1631 VSS.n1630 585
R1193 VSS.n1629 VSS.n1628 585
R1194 VSS.n1627 VSS.n1626 585
R1195 VSS.n1625 VSS.n1624 585
R1196 VSS.n1623 VSS.n1622 585
R1197 VSS.n1621 VSS.n903 585
R1198 VSS.n1621 VSS.n1620 585
R1199 VSS.n1597 VSS.n904 585
R1200 VSS.n905 VSS.n904 585
R1201 VSS.n1598 VSS.n911 585
R1202 VSS.n1612 VSS.n911 585
R1203 VSS.n1600 VSS.n918 585
R1204 VSS.n918 VSS.n910 585
R1205 VSS.n1603 VSS.n1602 585
R1206 VSS.n1605 VSS.n1603 585
R1207 VSS.n1596 VSS.n917 585
R1208 VSS.n1579 VSS.n917 585
R1209 VSS.n1595 VSS.n1594 585
R1210 VSS.n1594 VSS.n1593 585
R1211 VSS.n920 VSS.n919 585
R1212 VSS.n927 VSS.n920 585
R1213 VSS.n1562 VSS.n926 585
R1214 VSS.n1587 VSS.n926 585
R1215 VSS.n1564 VSS.n1563 585
R1216 VSS.n1565 VSS.n1564 585
R1217 VSS.n1561 VSS.n1044 585
R1218 VSS.n1050 VSS.n1044 585
R1219 VSS.n1560 VSS.n1559 585
R1220 VSS.n1559 VSS.n1558 585
R1221 VSS.n424 VSS.n217 394
R1222 VSS.n428 VSS.n217 394
R1223 VSS.n428 VSS.n211 394
R1224 VSS.n2199 VSS.n211 394
R1225 VSS.n2199 VSS.n209 394
R1226 VSS.n2203 VSS.n209 394
R1227 VSS.n2203 VSS.n204 394
R1228 VSS.n2212 VSS.n204 394
R1229 VSS.n2212 VSS.n202 394
R1230 VSS.n2216 VSS.n202 394
R1231 VSS.n2216 VSS.n197 394
R1232 VSS.n2225 VSS.n197 394
R1233 VSS.n2225 VSS.n195 394
R1234 VSS.n2229 VSS.n195 394
R1235 VSS.n2229 VSS.n190 394
R1236 VSS.n2238 VSS.n190 394
R1237 VSS.n2238 VSS.n188 394
R1238 VSS.n2242 VSS.n188 394
R1239 VSS.n2242 VSS.n183 394
R1240 VSS.n2251 VSS.n183 394
R1241 VSS.n2251 VSS.n181 394
R1242 VSS.n2255 VSS.n181 394
R1243 VSS.n2255 VSS.n176 394
R1244 VSS.n2263 VSS.n176 394
R1245 VSS.n2263 VSS.n174 394
R1246 VSS.n2267 VSS.n174 394
R1247 VSS.n2267 VSS.n168 394
R1248 VSS.n2275 VSS.n168 394
R1249 VSS.n2275 VSS.n166 394
R1250 VSS.n2279 VSS.n166 394
R1251 VSS.n2279 VSS.n160 394
R1252 VSS.n2287 VSS.n160 394
R1253 VSS.n2287 VSS.n158 394
R1254 VSS.n2291 VSS.n158 394
R1255 VSS.n2291 VSS.n152 394
R1256 VSS.n2299 VSS.n152 394
R1257 VSS.n2299 VSS.n150 394
R1258 VSS.n2303 VSS.n150 394
R1259 VSS.n2303 VSS.n144 394
R1260 VSS.n2311 VSS.n144 394
R1261 VSS.n2311 VSS.n142 394
R1262 VSS.n2315 VSS.n142 394
R1263 VSS.n2315 VSS.n136 394
R1264 VSS.n2323 VSS.n136 394
R1265 VSS.n2323 VSS.n134 394
R1266 VSS.n2327 VSS.n134 394
R1267 VSS.n2327 VSS.n128 394
R1268 VSS.n2335 VSS.n128 394
R1269 VSS.n2335 VSS.n126 394
R1270 VSS.n2339 VSS.n126 394
R1271 VSS.n2339 VSS.n120 394
R1272 VSS.n2347 VSS.n120 394
R1273 VSS.n2347 VSS.n118 394
R1274 VSS.n2351 VSS.n118 394
R1275 VSS.n2351 VSS.n112 394
R1276 VSS.n2359 VSS.n112 394
R1277 VSS.n2359 VSS.n110 394
R1278 VSS.n2363 VSS.n110 394
R1279 VSS.n2363 VSS.n103 394
R1280 VSS.n2398 VSS.n103 394
R1281 VSS.n2398 VSS.n101 394
R1282 VSS.n243 VSS.n219 394
R1283 VSS.n247 VSS.n241 394
R1284 VSS.n251 VSS.n249 394
R1285 VSS.n255 VSS.n239 394
R1286 VSS.n259 VSS.n257 394
R1287 VSS.n263 VSS.n237 394
R1288 VSS.n267 VSS.n265 394
R1289 VSS.n271 VSS.n235 394
R1290 VSS.n275 VSS.n273 394
R1291 VSS.n279 VSS.n233 394
R1292 VSS.n283 VSS.n281 394
R1293 VSS.n390 VSS.n229 394
R1294 VSS.n394 VSS.n392 394
R1295 VSS.n398 VSS.n227 394
R1296 VSS.n402 VSS.n400 394
R1297 VSS.n406 VSS.n225 394
R1298 VSS.n410 VSS.n408 394
R1299 VSS.n414 VSS.n223 394
R1300 VSS.n418 VSS.n416 394
R1301 VSS.n422 VSS.n215 394
R1302 VSS.n430 VSS.n215 394
R1303 VSS.n430 VSS.n213 394
R1304 VSS.n434 VSS.n213 394
R1305 VSS.n434 VSS.n208 394
R1306 VSS.n2205 VSS.n208 394
R1307 VSS.n2205 VSS.n206 394
R1308 VSS.n2209 VSS.n206 394
R1309 VSS.n2209 VSS.n201 394
R1310 VSS.n2218 VSS.n201 394
R1311 VSS.n2218 VSS.n199 394
R1312 VSS.n2222 VSS.n199 394
R1313 VSS.n2222 VSS.n194 394
R1314 VSS.n2231 VSS.n194 394
R1315 VSS.n2231 VSS.n192 394
R1316 VSS.n2235 VSS.n192 394
R1317 VSS.n2235 VSS.n187 394
R1318 VSS.n2244 VSS.n187 394
R1319 VSS.n2244 VSS.n185 394
R1320 VSS.n2248 VSS.n185 394
R1321 VSS.n2248 VSS.n180 394
R1322 VSS.n2257 VSS.n180 394
R1323 VSS.n2257 VSS.n178 394
R1324 VSS.n2261 VSS.n178 394
R1325 VSS.n2261 VSS.n172 394
R1326 VSS.n2269 VSS.n172 394
R1327 VSS.n2269 VSS.n170 394
R1328 VSS.n2273 VSS.n170 394
R1329 VSS.n2273 VSS.n164 394
R1330 VSS.n2281 VSS.n164 394
R1331 VSS.n2281 VSS.n162 394
R1332 VSS.n2285 VSS.n162 394
R1333 VSS.n2285 VSS.n156 394
R1334 VSS.n2293 VSS.n156 394
R1335 VSS.n2293 VSS.n154 394
R1336 VSS.n2297 VSS.n154 394
R1337 VSS.n2297 VSS.n147 394
R1338 VSS.n2305 VSS.n147 394
R1339 VSS.n2305 VSS.n145 394
R1340 VSS.n2309 VSS.n145 394
R1341 VSS.n2309 VSS.n139 394
R1342 VSS.n2317 VSS.n139 394
R1343 VSS.n2317 VSS.n137 394
R1344 VSS.n2321 VSS.n137 394
R1345 VSS.n2321 VSS.n131 394
R1346 VSS.n2329 VSS.n131 394
R1347 VSS.n2329 VSS.n129 394
R1348 VSS.n2333 VSS.n129 394
R1349 VSS.n2333 VSS.n123 394
R1350 VSS.n2341 VSS.n123 394
R1351 VSS.n2341 VSS.n121 394
R1352 VSS.n2345 VSS.n121 394
R1353 VSS.n2345 VSS.n115 394
R1354 VSS.n2353 VSS.n115 394
R1355 VSS.n2353 VSS.n113 394
R1356 VSS.n2357 VSS.n113 394
R1357 VSS.n2357 VSS.n108 394
R1358 VSS.n2365 VSS.n108 394
R1359 VSS.n2365 VSS.n105 394
R1360 VSS.n2396 VSS.n105 394
R1361 VSS.n2396 VSS.n106 394
R1362 VSS.n100 VSS.n99 394
R1363 VSS.n2443 VSS.n99 394
R1364 VSS.n2441 VSS.n2440 394
R1365 VSS.n2437 VSS.n2436 394
R1366 VSS.n2433 VSS.n2432 394
R1367 VSS.n2429 VSS.n2428 394
R1368 VSS.n2425 VSS.n2424 394
R1369 VSS.n2421 VSS.n2420 394
R1370 VSS.n2417 VSS.n2416 394
R1371 VSS.n2413 VSS.n2412 394
R1372 VSS.n2403 VSS.n2402 394
R1373 VSS.n2406 VSS.n79 394
R1374 VSS.n2452 VSS.n78 394
R1375 VSS.n2370 VSS.n2369 394
R1376 VSS.n2374 VSS.n2373 394
R1377 VSS.n2378 VSS.n2377 394
R1378 VSS.n2382 VSS.n2381 394
R1379 VSS.n2386 VSS.n2385 394
R1380 VSS.n2390 VSS.n2389 394
R1381 VSS.n1750 VSS.n876 394
R1382 VSS.n1750 VSS.n874 394
R1383 VSS.n1754 VSS.n874 394
R1384 VSS.n1754 VSS.n847 394
R1385 VSS.n1827 VSS.n847 394
R1386 VSS.n1827 VSS.n848 394
R1387 VSS.n848 VSS.n841 394
R1388 VSS.n1822 VSS.n841 394
R1389 VSS.n1822 VSS.n1821 394
R1390 VSS.n1821 VSS.n851 394
R1391 VSS.n1817 VSS.n851 394
R1392 VSS.n1736 VSS.n1686 394
R1393 VSS.n1732 VSS.n1731 394
R1394 VSS.n1728 VSS.n1727 394
R1395 VSS.n1724 VSS.n1723 394
R1396 VSS.n1720 VSS.n1719 394
R1397 VSS.n1716 VSS.n1715 394
R1398 VSS.n1712 VSS.n1711 394
R1399 VSS.n1708 VSS.n1707 394
R1400 VSS.n1704 VSS.n1703 394
R1401 VSS.n1700 VSS.n1699 394
R1402 VSS.n1696 VSS.n1695 394
R1403 VSS.n1691 VSS.n878 394
R1404 VSS.n878 VSS.n871 394
R1405 VSS.n1756 VSS.n871 394
R1406 VSS.n1758 VSS.n1756 394
R1407 VSS.n1758 VSS.n846 394
R1408 VSS.n1761 VSS.n846 394
R1409 VSS.n1761 VSS.n839 394
R1410 VSS.n1764 VSS.n839 394
R1411 VSS.n1764 VSS.n852 394
R1412 VSS.n853 VSS.n852 394
R1413 VSS.n854 VSS.n853 394
R1414 VSS.n1813 VSS.n1811 394
R1415 VSS.n1811 VSS.n1810 394
R1416 VSS.n1807 VSS.n1806 394
R1417 VSS.n1804 VSS.n861 394
R1418 VSS.n1800 VSS.n1798 394
R1419 VSS.n1796 VSS.n863 394
R1420 VSS.n1790 VSS.n1788 394
R1421 VSS.n1786 VSS.n866 394
R1422 VSS.n1782 VSS.n1780 394
R1423 VSS.n1778 VSS.n868 394
R1424 VSS.n1774 VSS.n1772 394
R1425 VSS.n1453 VSS.n1393 394
R1426 VSS.n1453 VSS.n1145 394
R1427 VSS.n1461 VSS.n1145 394
R1428 VSS.n1461 VSS.n1143 394
R1429 VSS.n1465 VSS.n1143 394
R1430 VSS.n1465 VSS.n1136 394
R1431 VSS.n1478 VSS.n1136 394
R1432 VSS.n1478 VSS.n1133 394
R1433 VSS.n1483 VSS.n1133 394
R1434 VSS.n1483 VSS.n1134 394
R1435 VSS.n1134 VSS.n1119 394
R1436 VSS.n1449 VSS.n1448 394
R1437 VSS.n1446 VSS.n1395 394
R1438 VSS.n1442 VSS.n1441 394
R1439 VSS.n1439 VSS.n1398 394
R1440 VSS.n1435 VSS.n1434 394
R1441 VSS.n1432 VSS.n1401 394
R1442 VSS.n1428 VSS.n1427 394
R1443 VSS.n1425 VSS.n1404 394
R1444 VSS.n1421 VSS.n1420 394
R1445 VSS.n1418 VSS.n1407 394
R1446 VSS.n1414 VSS.n1413 394
R1447 VSS.n1455 VSS.n1149 394
R1448 VSS.n1455 VSS.n1147 394
R1449 VSS.n1459 VSS.n1147 394
R1450 VSS.n1459 VSS.n1141 394
R1451 VSS.n1467 VSS.n1141 394
R1452 VSS.n1467 VSS.n1138 394
R1453 VSS.n1476 VSS.n1138 394
R1454 VSS.n1476 VSS.n1139 394
R1455 VSS.n1139 VSS.n1131 394
R1456 VSS.n1131 VSS.n1122 394
R1457 VSS.n1494 VSS.n1122 394
R1458 VSS.n1118 VSS.n1117 394
R1459 VSS.n1533 VSS.n1117 394
R1460 VSS.n1531 VSS.n1530 394
R1461 VSS.n1527 VSS.n1526 394
R1462 VSS.n1523 VSS.n1522 394
R1463 VSS.n1519 VSS.n1518 394
R1464 VSS.n1515 VSS.n1514 394
R1465 VSS.n1511 VSS.n1510 394
R1466 VSS.n1507 VSS.n1506 394
R1467 VSS.n1503 VSS.n1502 394
R1468 VSS.n1499 VSS.n1498 394
R1469 VSS.n2092 VSS.n648 394
R1470 VSS.n2088 VSS.n648 394
R1471 VSS.n2088 VSS.n651 394
R1472 VSS.n2084 VSS.n651 394
R1473 VSS.n2084 VSS.n653 394
R1474 VSS.n2080 VSS.n653 394
R1475 VSS.n2080 VSS.n655 394
R1476 VSS.n2076 VSS.n655 394
R1477 VSS.n2076 VSS.n657 394
R1478 VSS.n2072 VSS.n657 394
R1479 VSS.n2072 VSS.n659 394
R1480 VSS.n2068 VSS.n659 394
R1481 VSS.n2068 VSS.n661 394
R1482 VSS.n2064 VSS.n661 394
R1483 VSS.n2064 VSS.n663 394
R1484 VSS.n2060 VSS.n663 394
R1485 VSS.n2060 VSS.n665 394
R1486 VSS.n1042 VSS.n665 394
R1487 VSS.n1042 VSS.n1041 394
R1488 VSS.n1041 VSS.n1038 394
R1489 VSS.n1038 VSS.n770 394
R1490 VSS.n2049 VSS.n770 394
R1491 VSS.n2049 VSS.n771 394
R1492 VSS.n2045 VSS.n771 394
R1493 VSS.n2045 VSS.n773 394
R1494 VSS.n2041 VSS.n773 394
R1495 VSS.n2041 VSS.n776 394
R1496 VSS.n2037 VSS.n776 394
R1497 VSS.n2037 VSS.n778 394
R1498 VSS.n2033 VSS.n778 394
R1499 VSS.n2033 VSS.n780 394
R1500 VSS.n2029 VSS.n780 394
R1501 VSS.n2029 VSS.n782 394
R1502 VSS.n2025 VSS.n782 394
R1503 VSS.n2025 VSS.n784 394
R1504 VSS.n2021 VSS.n784 394
R1505 VSS.n2021 VSS.n786 394
R1506 VSS.n2017 VSS.n786 394
R1507 VSS.n1194 VSS.n1193 394
R1508 VSS.n1198 VSS.n1197 394
R1509 VSS.n1202 VSS.n1201 394
R1510 VSS.n1206 VSS.n1205 394
R1511 VSS.n1210 VSS.n1209 394
R1512 VSS.n1214 VSS.n1213 394
R1513 VSS.n1218 VSS.n1217 394
R1514 VSS.n1222 VSS.n1221 394
R1515 VSS.n1226 VSS.n1225 394
R1516 VSS.n1230 VSS.n1229 394
R1517 VSS.n1234 VSS.n1233 394
R1518 VSS.n1238 VSS.n1237 394
R1519 VSS.n1242 VSS.n1241 394
R1520 VSS.n1246 VSS.n1245 394
R1521 VSS.n1250 VSS.n1249 394
R1522 VSS.n1254 VSS.n1253 394
R1523 VSS.n1258 VSS.n1257 394
R1524 VSS.n1262 VSS.n1261 394
R1525 VSS.n1266 VSS.n1265 394
R1526 VSS.n1270 VSS.n1269 394
R1527 VSS.n1274 VSS.n1273 394
R1528 VSS.n1278 VSS.n1277 394
R1529 VSS.n1282 VSS.n1281 394
R1530 VSS.n1286 VSS.n1285 394
R1531 VSS.n1290 VSS.n1289 394
R1532 VSS.n1294 VSS.n1293 394
R1533 VSS.n1298 VSS.n1297 394
R1534 VSS.n1302 VSS.n1301 394
R1535 VSS.n1306 VSS.n1305 394
R1536 VSS.n1310 VSS.n1309 394
R1537 VSS.n1314 VSS.n1313 394
R1538 VSS.n1318 VSS.n1317 394
R1539 VSS.n1322 VSS.n1321 394
R1540 VSS.n1326 VSS.n1325 394
R1541 VSS.n1330 VSS.n1329 394
R1542 VSS.n1334 VSS.n1333 394
R1543 VSS.n1338 VSS.n1337 394
R1544 VSS.n1342 VSS.n1341 394
R1545 VSS.n1346 VSS.n1345 394
R1546 VSS.n1350 VSS.n1349 394
R1547 VSS.n1354 VSS.n1353 394
R1548 VSS.n1358 VSS.n1357 394
R1549 VSS.n1362 VSS.n1361 394
R1550 VSS.n1366 VSS.n1365 394
R1551 VSS.n1370 VSS.n1191 394
R1552 VSS.n1374 VSS.n1155 394
R1553 VSS.n1391 VSS.n1153 394
R1554 VSS.n1387 VSS.n1153 394
R1555 VSS.n1387 VSS.n1384 394
R1556 VSS.n1384 VSS.n1383 394
R1557 VSS.n1383 VSS.n1378 394
R1558 VSS.n1378 VSS.n1128 394
R1559 VSS.n1486 VSS.n1128 394
R1560 VSS.n1486 VSS.n1124 394
R1561 VSS.n1491 VSS.n1124 394
R1562 VSS.n1491 VSS.n1126 394
R1563 VSS.n1126 VSS.n1105 394
R1564 VSS.n1543 VSS.n1105 394
R1565 VSS.n1543 VSS.n1102 394
R1566 VSS.n1548 VSS.n1102 394
R1567 VSS.n1548 VSS.n1103 394
R1568 VSS.n1103 VSS.n1034 394
R1569 VSS.n1567 VSS.n1034 394
R1570 VSS.n1567 VSS.n928 394
R1571 VSS.n1585 VSS.n928 394
R1572 VSS.n1585 VSS.n929 394
R1573 VSS.n1581 VSS.n929 394
R1574 VSS.n1581 VSS.n1578 394
R1575 VSS.n1578 VSS.n909 394
R1576 VSS.n1614 VSS.n909 394
R1577 VSS.n1614 VSS.n907 394
R1578 VSS.n1618 VSS.n907 394
R1579 VSS.n1618 VSS.n887 394
R1580 VSS.n1669 VSS.n887 394
R1581 VSS.n1669 VSS.n885 394
R1582 VSS.n1673 VSS.n885 394
R1583 VSS.n1673 VSS.n883 394
R1584 VSS.n1740 VSS.n883 394
R1585 VSS.n1740 VSS.n880 394
R1586 VSS.n1747 VSS.n880 394
R1587 VSS.n1747 VSS.n881 394
R1588 VSS.n1743 VSS.n881 394
R1589 VSS.n1743 VSS.n844 394
R1590 VSS.n1830 VSS.n844 394
R1591 VSS.n2013 VSS.n799 394
R1592 VSS.n2009 VSS.n799 394
R1593 VSS.n2007 VSS.n2006 394
R1594 VSS.n2003 VSS.n2002 394
R1595 VSS.n1999 VSS.n1998 394
R1596 VSS.n1995 VSS.n1994 394
R1597 VSS.n1991 VSS.n1990 394
R1598 VSS.n1987 VSS.n1986 394
R1599 VSS.n1983 VSS.n1982 394
R1600 VSS.n1979 VSS.n798 394
R1601 VSS.n1976 VSS.n798 394
R1602 VSS.n1973 VSS.n801 394
R1603 VSS.n1969 VSS.n1968 394
R1604 VSS.n1965 VSS.n1964 394
R1605 VSS.n1961 VSS.n1960 394
R1606 VSS.n1957 VSS.n1956 394
R1607 VSS.n1953 VSS.n1952 394
R1608 VSS.n1949 VSS.n1948 394
R1609 VSS.n1945 VSS.n1944 394
R1610 VSS.n1941 VSS.n1940 394
R1611 VSS.n1937 VSS.n1936 394
R1612 VSS.n1933 VSS.n1932 394
R1613 VSS.n1929 VSS.n1928 394
R1614 VSS.n1921 VSS.n1920 394
R1615 VSS.n1917 VSS.n1916 394
R1616 VSS.n1913 VSS.n1912 394
R1617 VSS.n1909 VSS.n1908 394
R1618 VSS.n1905 VSS.n1904 394
R1619 VSS.n1901 VSS.n1900 394
R1620 VSS.n1897 VSS.n1896 394
R1621 VSS.n1893 VSS.n1892 394
R1622 VSS.n1889 VSS.n1888 394
R1623 VSS.n1885 VSS.n1884 394
R1624 VSS.n1881 VSS.n1880 394
R1625 VSS.n1873 VSS.n1872 394
R1626 VSS.n1869 VSS.n1868 394
R1627 VSS.n1865 VSS.n1864 394
R1628 VSS.n1861 VSS.n1860 394
R1629 VSS.n1857 VSS.n1856 394
R1630 VSS.n1853 VSS.n1852 394
R1631 VSS.n1849 VSS.n1848 394
R1632 VSS.n1845 VSS.n1844 394
R1633 VSS.n1841 VSS.n1840 394
R1634 VSS.n1837 VSS.n1836 394
R1635 VSS.n1833 VSS.n838 394
R1636 VSS.n543 VSS.n538 394
R1637 VSS.n547 VSS.n545 394
R1638 VSS.n553 VSS.n536 394
R1639 VSS.n557 VSS.n536 394
R1640 VSS.n557 VSS.n530 394
R1641 VSS.n566 VSS.n530 394
R1642 VSS.n566 VSS.n528 394
R1643 VSS.n570 VSS.n528 394
R1644 VSS.n570 VSS.n438 394
R1645 VSS.n2194 VSS.n438 394
R1646 VSS.n2194 VSS.n439 394
R1647 VSS.n2190 VSS.n439 394
R1648 VSS.n2190 VSS.n442 394
R1649 VSS.n2186 VSS.n442 394
R1650 VSS.n2186 VSS.n447 394
R1651 VSS.n2182 VSS.n447 394
R1652 VSS.n2182 VSS.n449 394
R1653 VSS.n2178 VSS.n449 394
R1654 VSS.n2178 VSS.n454 394
R1655 VSS.n2174 VSS.n454 394
R1656 VSS.n2174 VSS.n456 394
R1657 VSS.n2170 VSS.n456 394
R1658 VSS.n2170 VSS.n461 394
R1659 VSS.n2166 VSS.n461 394
R1660 VSS.n2166 VSS.n463 394
R1661 VSS.n2162 VSS.n463 394
R1662 VSS.n2162 VSS.n468 394
R1663 VSS.n2158 VSS.n468 394
R1664 VSS.n2158 VSS.n470 394
R1665 VSS.n2154 VSS.n470 394
R1666 VSS.n2154 VSS.n475 394
R1667 VSS.n2150 VSS.n475 394
R1668 VSS.n2150 VSS.n477 394
R1669 VSS.n2146 VSS.n477 394
R1670 VSS.n2146 VSS.n482 394
R1671 VSS.n2142 VSS.n482 394
R1672 VSS.n2142 VSS.n484 394
R1673 VSS.n2138 VSS.n484 394
R1674 VSS.n2138 VSS.n489 394
R1675 VSS.n2134 VSS.n489 394
R1676 VSS.n2134 VSS.n491 394
R1677 VSS.n2130 VSS.n491 394
R1678 VSS.n2130 VSS.n496 394
R1679 VSS.n2126 VSS.n496 394
R1680 VSS.n2126 VSS.n498 394
R1681 VSS.n2122 VSS.n498 394
R1682 VSS.n2122 VSS.n503 394
R1683 VSS.n2118 VSS.n503 394
R1684 VSS.n2118 VSS.n505 394
R1685 VSS.n2114 VSS.n505 394
R1686 VSS.n2114 VSS.n510 394
R1687 VSS.n2110 VSS.n510 394
R1688 VSS.n2110 VSS.n512 394
R1689 VSS.n2106 VSS.n512 394
R1690 VSS.n2106 VSS.n517 394
R1691 VSS.n2098 VSS.n521 394
R1692 VSS.n522 VSS.n521 394
R1693 VSS.n551 VSS.n534 394
R1694 VSS.n559 VSS.n534 394
R1695 VSS.n559 VSS.n532 394
R1696 VSS.n564 VSS.n532 394
R1697 VSS.n564 VSS.n526 394
R1698 VSS.n572 VSS.n526 394
R1699 VSS.n573 VSS.n572 394
R1700 VSS.n573 VSS.n436 394
R1701 VSS.n576 VSS.n436 394
R1702 VSS.n576 VSS.n443 394
R1703 VSS.n444 VSS.n443 394
R1704 VSS.n445 VSS.n444 394
R1705 VSS.n581 VSS.n445 394
R1706 VSS.n581 VSS.n450 394
R1707 VSS.n451 VSS.n450 394
R1708 VSS.n452 VSS.n451 394
R1709 VSS.n586 VSS.n452 394
R1710 VSS.n586 VSS.n457 394
R1711 VSS.n458 VSS.n457 394
R1712 VSS.n459 VSS.n458 394
R1713 VSS.n591 VSS.n459 394
R1714 VSS.n591 VSS.n464 394
R1715 VSS.n465 VSS.n464 394
R1716 VSS.n466 VSS.n465 394
R1717 VSS.n596 VSS.n466 394
R1718 VSS.n596 VSS.n471 394
R1719 VSS.n599 VSS.n471 394
R1720 VSS.n599 VSS.n473 394
R1721 VSS.n602 VSS.n473 394
R1722 VSS.n602 VSS.n478 394
R1723 VSS.n479 VSS.n478 394
R1724 VSS.n480 VSS.n479 394
R1725 VSS.n607 VSS.n480 394
R1726 VSS.n607 VSS.n485 394
R1727 VSS.n486 VSS.n485 394
R1728 VSS.n487 VSS.n486 394
R1729 VSS.n612 VSS.n487 394
R1730 VSS.n612 VSS.n492 394
R1731 VSS.n493 VSS.n492 394
R1732 VSS.n494 VSS.n493 394
R1733 VSS.n617 VSS.n494 394
R1734 VSS.n617 VSS.n499 394
R1735 VSS.n500 VSS.n499 394
R1736 VSS.n501 VSS.n500 394
R1737 VSS.n622 VSS.n501 394
R1738 VSS.n622 VSS.n506 394
R1739 VSS.n507 VSS.n506 394
R1740 VSS.n508 VSS.n507 394
R1741 VSS.n627 VSS.n508 394
R1742 VSS.n627 VSS.n513 394
R1743 VSS.n514 VSS.n513 394
R1744 VSS.n515 VSS.n514 394
R1745 VSS.n523 VSS.n515 394
R1746 VSS.n1557 VSS.n1051 394
R1747 VSS.n1051 VSS.n924 394
R1748 VSS.n1588 VSS.n924 394
R1749 VSS.n1588 VSS.n922 394
R1750 VSS.n1592 VSS.n922 394
R1751 VSS.n1592 VSS.n915 394
R1752 VSS.n1606 VSS.n915 394
R1753 VSS.n1606 VSS.n912 394
R1754 VSS.n1611 VSS.n912 394
R1755 VSS.n1611 VSS.n913 394
R1756 VSS.n913 VSS.n901 394
R1757 VSS.n900 VSS.n899 394
R1758 VSS.n1660 VSS.n899 394
R1759 VSS.n1658 VSS.n1657 394
R1760 VSS.n1654 VSS.n1653 394
R1761 VSS.n1650 VSS.n1649 394
R1762 VSS.n1646 VSS.n1645 394
R1763 VSS.n1642 VSS.n1641 394
R1764 VSS.n1638 VSS.n1637 394
R1765 VSS.n1634 VSS.n1633 394
R1766 VSS.n1630 VSS.n1629 394
R1767 VSS.n1626 VSS.n1625 394
R1768 VSS.n1559 VSS.n1044 394
R1769 VSS.n1564 VSS.n1044 394
R1770 VSS.n1564 VSS.n926 394
R1771 VSS.n926 VSS.n920 394
R1772 VSS.n1594 VSS.n920 394
R1773 VSS.n1594 VSS.n917 394
R1774 VSS.n1603 VSS.n917 394
R1775 VSS.n1603 VSS.n918 394
R1776 VSS.n918 VSS.n911 394
R1777 VSS.n911 VSS.n904 394
R1778 VSS.n1621 VSS.n904 394
R1779 VSS.n1552 VSS.n1053 394
R1780 VSS.n1066 VSS.n1065 394
R1781 VSS.n1070 VSS.n1069 394
R1782 VSS.n1074 VSS.n1073 394
R1783 VSS.n1078 VSS.n1077 394
R1784 VSS.n1082 VSS.n1081 394
R1785 VSS.n1086 VSS.n1085 394
R1786 VSS.n1090 VSS.n1089 394
R1787 VSS.n1094 VSS.n1093 394
R1788 VSS.n1096 VSS.n1063 394
R1789 VSS.n1100 VSS.n1046 394
R1790 VSS.n2155 VSS.n474 328.791
R1791 VSS.n2149 VSS.n474 328.791
R1792 VSS.n2149 VSS.n2148 328.791
R1793 VSS.n2148 VSS.n2147 328.791
R1794 VSS.n2147 VSS.n481 328.791
R1795 VSS.n2141 VSS.n481 328.791
R1796 VSS.n2141 VSS.n2140 328.791
R1797 VSS.n2140 VSS.n2139 328.791
R1798 VSS.n2139 VSS.n488 328.791
R1799 VSS.n2133 VSS.n488 328.791
R1800 VSS.n2133 VSS.n2132 328.791
R1801 VSS.n2132 VSS.n2131 328.791
R1802 VSS.n2131 VSS.n495 328.791
R1803 VSS.n2125 VSS.n495 328.791
R1804 VSS.n2125 VSS.n2124 328.791
R1805 VSS.n2124 VSS.n2123 328.791
R1806 VSS.n2123 VSS.n502 328.791
R1807 VSS.n2117 VSS.n502 328.791
R1808 VSS.n2117 VSS.n2116 328.791
R1809 VSS.n2116 VSS.n2115 328.791
R1810 VSS.n2115 VSS.n509 328.791
R1811 VSS.n2109 VSS.n509 328.791
R1812 VSS.n2109 VSS.n2108 328.791
R1813 VSS.n2108 VSS.n2107 328.791
R1814 VSS.n2107 VSS.n516 328.791
R1815 VSS.n71 VSS.n70 325.69
R1816 VSS.n16 VSS.n11 325.69
R1817 VSS.n1237 VSS.n1157 269.089
R1818 VSS.n1234 VSS.n1157 269.089
R1819 VSS.n2450 VSS.n98 261
R1820 VSS.n758 VSS.t81 259.341
R1821 VSS.n675 VSS.t35 259.341
R1822 VSS.n1021 VSS.t41 259.341
R1823 VSS.n938 VSS.t44 259.341
R1824 VSS.n757 VSS.t84 258.99
R1825 VSS.n756 VSS.t68 258.99
R1826 VSS.n755 VSS.t50 258.99
R1827 VSS.n668 VSS.t101 258.99
R1828 VSS.n669 VSS.t89 258.99
R1829 VSS.n672 VSS.t93 258.99
R1830 VSS.n673 VSS.t74 258.99
R1831 VSS.n674 VSS.t53 258.99
R1832 VSS.n1020 VSS.t91 258.99
R1833 VSS.n1019 VSS.t70 258.99
R1834 VSS.n1018 VSS.t72 258.99
R1835 VSS.n931 VSS.t76 258.99
R1836 VSS.n932 VSS.t78 258.99
R1837 VSS.n935 VSS.t103 258.99
R1838 VSS.n936 VSS.t33 258.99
R1839 VSS.n937 VSS.t38 258.99
R1840 VSS.n750 VSS.n720 253.042
R1841 VSS.n690 VSS.n689 253.042
R1842 VSS.n1016 VSS.n1015 253.042
R1843 VSS.n952 VSS.n949 253.042
R1844 VSS.n546 VSS.n539 218.815
R1845 VSS.n544 VSS.n539 218.815
R1846 VSS.n2097 VSS.n2095 218.815
R1847 VSS.n2095 VSS.n635 218.815
R1848 VSS.n2015 VSS.n2014 218.815
R1849 VSS.n2015 VSS.n790 218.815
R1850 VSS.n2015 VSS.n791 218.815
R1851 VSS.n2015 VSS.n792 218.815
R1852 VSS.n2015 VSS.n793 218.815
R1853 VSS.n2015 VSS.n794 218.815
R1854 VSS.n2015 VSS.n795 218.815
R1855 VSS.n2015 VSS.n796 218.815
R1856 VSS.n2015 VSS.n797 218.815
R1857 VSS.n2094 VSS.n645 218.815
R1858 VSS.n2094 VSS.n644 218.815
R1859 VSS.n2094 VSS.n643 218.815
R1860 VSS.n2094 VSS.n642 218.815
R1861 VSS.n2094 VSS.n641 218.815
R1862 VSS.n2094 VSS.n640 218.815
R1863 VSS.n2094 VSS.n639 218.815
R1864 VSS.n2094 VSS.n638 218.815
R1865 VSS.n2094 VSS.n637 218.815
R1866 VSS.n2094 VSS.n636 218.815
R1867 VSS.n1540 VSS.n1539 218.815
R1868 VSS.n1540 VSS.n1107 218.815
R1869 VSS.n1540 VSS.n1108 218.815
R1870 VSS.n1540 VSS.n1109 218.815
R1871 VSS.n1540 VSS.n1110 218.815
R1872 VSS.n1540 VSS.n1111 218.815
R1873 VSS.n1540 VSS.n1112 218.815
R1874 VSS.n1540 VSS.n1113 218.815
R1875 VSS.n1540 VSS.n1114 218.815
R1876 VSS.n1540 VSS.n1115 218.815
R1877 VSS.n1540 VSS.n1116 218.815
R1878 VSS.n1412 VSS.n98 218.815
R1879 VSS.n1409 VSS.n98 218.815
R1880 VSS.n1419 VSS.n98 218.815
R1881 VSS.n1406 VSS.n98 218.815
R1882 VSS.n1426 VSS.n98 218.815
R1883 VSS.n1403 VSS.n98 218.815
R1884 VSS.n1433 VSS.n98 218.815
R1885 VSS.n1400 VSS.n98 218.815
R1886 VSS.n1440 VSS.n98 218.815
R1887 VSS.n1397 VSS.n98 218.815
R1888 VSS.n1447 VSS.n98 218.815
R1889 VSS.n1812 VSS.n855 218.815
R1890 VSS.n859 VSS.n855 218.815
R1891 VSS.n1805 VSS.n855 218.815
R1892 VSS.n1799 VSS.n855 218.815
R1893 VSS.n1797 VSS.n855 218.815
R1894 VSS.n1789 VSS.n855 218.815
R1895 VSS.n1787 VSS.n855 218.815
R1896 VSS.n1781 VSS.n855 218.815
R1897 VSS.n1779 VSS.n855 218.815
R1898 VSS.n1773 VSS.n855 218.815
R1899 VSS.n1771 VSS.n855 218.815
R1900 VSS.n1737 VSS.n1675 218.815
R1901 VSS.n1737 VSS.n1676 218.815
R1902 VSS.n1737 VSS.n1677 218.815
R1903 VSS.n1737 VSS.n1678 218.815
R1904 VSS.n1737 VSS.n1679 218.815
R1905 VSS.n1737 VSS.n1680 218.815
R1906 VSS.n1737 VSS.n1681 218.815
R1907 VSS.n1737 VSS.n1682 218.815
R1908 VSS.n1737 VSS.n1683 218.815
R1909 VSS.n1737 VSS.n1684 218.815
R1910 VSS.n1737 VSS.n1685 218.815
R1911 VSS.n2450 VSS.n2449 218.815
R1912 VSS.n2450 VSS.n81 218.815
R1913 VSS.n2450 VSS.n82 218.815
R1914 VSS.n2450 VSS.n83 218.815
R1915 VSS.n2450 VSS.n84 218.815
R1916 VSS.n2450 VSS.n85 218.815
R1917 VSS.n2450 VSS.n86 218.815
R1918 VSS.n2450 VSS.n87 218.815
R1919 VSS.n2450 VSS.n88 218.815
R1920 VSS.n2450 VSS.n89 218.815
R1921 VSS.n2450 VSS.n90 218.815
R1922 VSS.n2451 VSS.n2450 218.815
R1923 VSS.n2450 VSS.n91 218.815
R1924 VSS.n2450 VSS.n92 218.815
R1925 VSS.n2450 VSS.n93 218.815
R1926 VSS.n2450 VSS.n94 218.815
R1927 VSS.n2450 VSS.n95 218.815
R1928 VSS.n2450 VSS.n96 218.815
R1929 VSS.n2450 VSS.n97 218.815
R1930 VSS.n417 VSS.n220 218.815
R1931 VSS.n415 VSS.n220 218.815
R1932 VSS.n409 VSS.n220 218.815
R1933 VSS.n407 VSS.n220 218.815
R1934 VSS.n401 VSS.n220 218.815
R1935 VSS.n399 VSS.n220 218.815
R1936 VSS.n393 VSS.n220 218.815
R1937 VSS.n391 VSS.n220 218.815
R1938 VSS.n282 VSS.n220 218.815
R1939 VSS.n280 VSS.n220 218.815
R1940 VSS.n274 VSS.n220 218.815
R1941 VSS.n272 VSS.n220 218.815
R1942 VSS.n266 VSS.n220 218.815
R1943 VSS.n264 VSS.n220 218.815
R1944 VSS.n258 VSS.n220 218.815
R1945 VSS.n256 VSS.n220 218.815
R1946 VSS.n250 VSS.n220 218.815
R1947 VSS.n248 VSS.n220 218.815
R1948 VSS.n242 VSS.n220 218.815
R1949 VSS.n1975 VSS.n1974 218.815
R1950 VSS.n1974 VSS.n803 218.815
R1951 VSS.n1974 VSS.n804 218.815
R1952 VSS.n1974 VSS.n805 218.815
R1953 VSS.n1974 VSS.n806 218.815
R1954 VSS.n1974 VSS.n807 218.815
R1955 VSS.n1974 VSS.n808 218.815
R1956 VSS.n1974 VSS.n809 218.815
R1957 VSS.n1974 VSS.n810 218.815
R1958 VSS.n1974 VSS.n811 218.815
R1959 VSS.n1974 VSS.n812 218.815
R1960 VSS.n1974 VSS.n813 218.815
R1961 VSS.n1974 VSS.n814 218.815
R1962 VSS.n1974 VSS.n815 218.815
R1963 VSS.n1974 VSS.n816 218.815
R1964 VSS.n1974 VSS.n817 218.815
R1965 VSS.n1974 VSS.n818 218.815
R1966 VSS.n1974 VSS.n819 218.815
R1967 VSS.n1974 VSS.n820 218.815
R1968 VSS.n1974 VSS.n821 218.815
R1969 VSS.n1974 VSS.n822 218.815
R1970 VSS.n1974 VSS.n823 218.815
R1971 VSS.n1974 VSS.n824 218.815
R1972 VSS.n1974 VSS.n825 218.815
R1973 VSS.n1974 VSS.n826 218.815
R1974 VSS.n1974 VSS.n827 218.815
R1975 VSS.n1974 VSS.n828 218.815
R1976 VSS.n1974 VSS.n829 218.815
R1977 VSS.n1974 VSS.n830 218.815
R1978 VSS.n1974 VSS.n831 218.815
R1979 VSS.n1974 VSS.n832 218.815
R1980 VSS.n1974 VSS.n833 218.815
R1981 VSS.n1974 VSS.n834 218.815
R1982 VSS.n1974 VSS.n835 218.815
R1983 VSS.n1974 VSS.n836 218.815
R1984 VSS.n1974 VSS.n837 218.815
R1985 VSS.n1373 VSS.n1372 218.815
R1986 VSS.n1372 VSS.n1371 218.815
R1987 VSS.n1372 VSS.n1190 218.815
R1988 VSS.n1372 VSS.n1189 218.815
R1989 VSS.n1372 VSS.n1188 218.815
R1990 VSS.n1372 VSS.n1187 218.815
R1991 VSS.n1372 VSS.n1186 218.815
R1992 VSS.n1372 VSS.n1185 218.815
R1993 VSS.n1372 VSS.n1184 218.815
R1994 VSS.n1372 VSS.n1183 218.815
R1995 VSS.n1372 VSS.n1182 218.815
R1996 VSS.n1372 VSS.n1180 218.815
R1997 VSS.n1372 VSS.n1179 218.815
R1998 VSS.n1372 VSS.n1178 218.815
R1999 VSS.n1372 VSS.n1177 218.815
R2000 VSS.n1372 VSS.n1176 218.815
R2001 VSS.n1372 VSS.n1175 218.815
R2002 VSS.n1372 VSS.n1174 218.815
R2003 VSS.n1372 VSS.n1173 218.815
R2004 VSS.n1372 VSS.n1172 218.815
R2005 VSS.n1372 VSS.n1171 218.815
R2006 VSS.n1372 VSS.n1170 218.815
R2007 VSS.n1372 VSS.n1168 218.815
R2008 VSS.n1372 VSS.n1167 218.815
R2009 VSS.n1372 VSS.n1166 218.815
R2010 VSS.n1372 VSS.n1165 218.815
R2011 VSS.n1372 VSS.n1164 218.815
R2012 VSS.n1372 VSS.n1163 218.815
R2013 VSS.n1372 VSS.n1162 218.815
R2014 VSS.n1372 VSS.n1161 218.815
R2015 VSS.n1372 VSS.n1160 218.815
R2016 VSS.n1372 VSS.n1159 218.815
R2017 VSS.n1372 VSS.n1158 218.815
R2018 VSS.n1372 VSS.n1156 218.815
R2019 VSS.n1550 VSS.n1101 218.815
R2020 VSS.n1550 VSS.n1062 218.815
R2021 VSS.n1550 VSS.n1061 218.815
R2022 VSS.n1550 VSS.n1060 218.815
R2023 VSS.n1550 VSS.n1059 218.815
R2024 VSS.n1550 VSS.n1058 218.815
R2025 VSS.n1550 VSS.n1057 218.815
R2026 VSS.n1550 VSS.n1056 218.815
R2027 VSS.n1550 VSS.n1055 218.815
R2028 VSS.n1550 VSS.n1054 218.815
R2029 VSS.n1551 VSS.n1550 218.815
R2030 VSS.n1667 VSS.n1666 218.815
R2031 VSS.n1667 VSS.n889 218.815
R2032 VSS.n1667 VSS.n890 218.815
R2033 VSS.n1667 VSS.n891 218.815
R2034 VSS.n1667 VSS.n892 218.815
R2035 VSS.n1667 VSS.n893 218.815
R2036 VSS.n1667 VSS.n894 218.815
R2037 VSS.n1667 VSS.n895 218.815
R2038 VSS.n1667 VSS.n896 218.815
R2039 VSS.n1667 VSS.n897 218.815
R2040 VSS.n1667 VSS.n898 218.815
R2041 VSS.n1285 VSS.n1169 198.87
R2042 VSS.n1333 VSS.n1181 198.87
R2043 VSS.n1330 VSS.n1181 198.87
R2044 VSS.n1282 VSS.n1169 198.87
R2045 VSS.n1372 VSS.n1181 193.066
R2046 VSS.n1372 VSS.n1169 193.066
R2047 VSS.n552 VSS.n539 185.895
R2048 VSS.n320 VSS.n319 185
R2049 VSS.n320 VSS.n292 185
R2050 VSS.n322 VSS.n321 185
R2051 VSS.n321 VSS.n290 185
R2052 VSS.n304 VSS.n296 185
R2053 VSS.n304 VSS.n295 185
R2054 VSS.n305 VSS.n304 185
R2055 VSS.n382 VSS.n381 185
R2056 VSS.n381 VSS.n365 185
R2057 VSS.n380 VSS.n379 185
R2058 VSS.n380 VSS.n367 185
R2059 VSS.n359 VSS.n351 185
R2060 VSS.n359 VSS.n350 185
R2061 VSS.n360 VSS.n359 185
R2062 VSS.n70 VSS.n69 185
R2063 VSS.n47 VSS.n46 185
R2064 VSS.n64 VSS.n63 185
R2065 VSS.n58 VSS.n57 185
R2066 VSS.n58 VSS.n50 185
R2067 VSS.n30 VSS.n29 185
R2068 VSS.n29 VSS.n28 185
R2069 VSS.n16 VSS.n15 185
R2070 VSS.n18 VSS.n17 185
R2071 VSS.n20 VSS.n8 185
R2072 VSS.n751 VSS.n750 185
R2073 VSS.n749 VSS.n748 185
R2074 VSS.n724 VSS.n723 185
R2075 VSS.n743 VSS.n742 185
R2076 VSS.n741 VSS.n740 185
R2077 VSS.n728 VSS.n727 185
R2078 VSS.n735 VSS.n734 185
R2079 VSS.n733 VSS.n732 185
R2080 VSS.n691 VSS.n690 185
R2081 VSS.n685 VSS.n684 185
R2082 VSS.n697 VSS.n696 185
R2083 VSS.n699 VSS.n698 185
R2084 VSS.n681 VSS.n680 185
R2085 VSS.n706 VSS.n705 185
R2086 VSS.n708 VSS.n707 185
R2087 VSS.n710 VSS.n677 185
R2088 VSS.n994 VSS.n993 185
R2089 VSS.n999 VSS.n998 185
R2090 VSS.n1001 VSS.n1000 185
R2091 VSS.n990 VSS.n989 185
R2092 VSS.n1007 VSS.n1006 185
R2093 VSS.n1009 VSS.n1008 185
R2094 VSS.n986 VSS.n985 185
R2095 VSS.n1015 VSS.n1014 185
R2096 VSS.n974 VSS.n973 185
R2097 VSS.n942 VSS.n941 185
R2098 VSS.n968 VSS.n967 185
R2099 VSS.n966 VSS.n965 185
R2100 VSS.n946 VSS.n945 185
R2101 VSS.n960 VSS.n959 185
R2102 VSS.n958 VSS.n957 185
R2103 VSS.n950 VSS.n949 185
R2104 VSS.n731 VSS.t83 178.418
R2105 VSS.t37 VSS.n711 178.418
R2106 VSS.n995 VSS.t43 178.418
R2107 VSS.t45 VSS.n940 178.418
R2108 VSS.t88 VSS.n62 175.332
R2109 VSS.t98 VSS.n21 175.332
R2110 VSS.n2094 VSS.n2093 163.94
R2111 VSS.n2016 VSS.n2015 163.94
R2112 VSS.n1372 VSS.n1157 157.957
R2113 VSS.n242 VSS.n241 147.374
R2114 VSS.n249 VSS.n248 147.374
R2115 VSS.n250 VSS.n239 147.374
R2116 VSS.n257 VSS.n256 147.374
R2117 VSS.n258 VSS.n237 147.374
R2118 VSS.n265 VSS.n264 147.374
R2119 VSS.n266 VSS.n235 147.374
R2120 VSS.n273 VSS.n272 147.374
R2121 VSS.n274 VSS.n233 147.374
R2122 VSS.n281 VSS.n280 147.374
R2123 VSS.n282 VSS.n229 147.374
R2124 VSS.n392 VSS.n391 147.374
R2125 VSS.n393 VSS.n227 147.374
R2126 VSS.n400 VSS.n399 147.374
R2127 VSS.n401 VSS.n225 147.374
R2128 VSS.n408 VSS.n407 147.374
R2129 VSS.n409 VSS.n223 147.374
R2130 VSS.n416 VSS.n415 147.374
R2131 VSS.n417 VSS.n221 147.374
R2132 VSS.n2449 VSS.n2448 147.374
R2133 VSS.n2443 VSS.n81 147.374
R2134 VSS.n2440 VSS.n82 147.374
R2135 VSS.n2436 VSS.n83 147.374
R2136 VSS.n2432 VSS.n84 147.374
R2137 VSS.n2428 VSS.n85 147.374
R2138 VSS.n2424 VSS.n86 147.374
R2139 VSS.n2420 VSS.n87 147.374
R2140 VSS.n2416 VSS.n88 147.374
R2141 VSS.n2412 VSS.n89 147.374
R2142 VSS.n2403 VSS.n90 147.374
R2143 VSS.n2451 VSS.n79 147.374
R2144 VSS.n91 VSS.n78 147.374
R2145 VSS.n2370 VSS.n92 147.374
R2146 VSS.n2374 VSS.n93 147.374
R2147 VSS.n2378 VSS.n94 147.374
R2148 VSS.n2382 VSS.n95 147.374
R2149 VSS.n2386 VSS.n96 147.374
R2150 VSS.n2390 VSS.n97 147.374
R2151 VSS.n1732 VSS.n1685 147.374
R2152 VSS.n1728 VSS.n1684 147.374
R2153 VSS.n1724 VSS.n1683 147.374
R2154 VSS.n1720 VSS.n1682 147.374
R2155 VSS.n1716 VSS.n1681 147.374
R2156 VSS.n1712 VSS.n1680 147.374
R2157 VSS.n1708 VSS.n1679 147.374
R2158 VSS.n1704 VSS.n1678 147.374
R2159 VSS.n1700 VSS.n1677 147.374
R2160 VSS.n1696 VSS.n1676 147.374
R2161 VSS.n1692 VSS.n1675 147.374
R2162 VSS.n1812 VSS.n856 147.374
R2163 VSS.n1810 VSS.n859 147.374
R2164 VSS.n1806 VSS.n1805 147.374
R2165 VSS.n1799 VSS.n861 147.374
R2166 VSS.n1798 VSS.n1797 147.374
R2167 VSS.n1789 VSS.n863 147.374
R2168 VSS.n1788 VSS.n1787 147.374
R2169 VSS.n1781 VSS.n866 147.374
R2170 VSS.n1780 VSS.n1779 147.374
R2171 VSS.n1773 VSS.n868 147.374
R2172 VSS.n1772 VSS.n1771 147.374
R2173 VSS.n1447 VSS.n1446 147.374
R2174 VSS.n1442 VSS.n1397 147.374
R2175 VSS.n1440 VSS.n1439 147.374
R2176 VSS.n1435 VSS.n1400 147.374
R2177 VSS.n1433 VSS.n1432 147.374
R2178 VSS.n1428 VSS.n1403 147.374
R2179 VSS.n1426 VSS.n1425 147.374
R2180 VSS.n1421 VSS.n1406 147.374
R2181 VSS.n1419 VSS.n1418 147.374
R2182 VSS.n1414 VSS.n1409 147.374
R2183 VSS.n1412 VSS.n1411 147.374
R2184 VSS.n1539 VSS.n1538 147.374
R2185 VSS.n1533 VSS.n1107 147.374
R2186 VSS.n1530 VSS.n1108 147.374
R2187 VSS.n1526 VSS.n1109 147.374
R2188 VSS.n1522 VSS.n1110 147.374
R2189 VSS.n1518 VSS.n1111 147.374
R2190 VSS.n1514 VSS.n1112 147.374
R2191 VSS.n1510 VSS.n1113 147.374
R2192 VSS.n1506 VSS.n1114 147.374
R2193 VSS.n1502 VSS.n1115 147.374
R2194 VSS.n1498 VSS.n1116 147.374
R2195 VSS.n1193 VSS.n636 147.374
R2196 VSS.n1197 VSS.n637 147.374
R2197 VSS.n1201 VSS.n638 147.374
R2198 VSS.n1205 VSS.n639 147.374
R2199 VSS.n1209 VSS.n640 147.374
R2200 VSS.n1213 VSS.n641 147.374
R2201 VSS.n1217 VSS.n642 147.374
R2202 VSS.n1221 VSS.n643 147.374
R2203 VSS.n1225 VSS.n644 147.374
R2204 VSS.n1229 VSS.n645 147.374
R2205 VSS.n1233 VSS.n1156 147.374
R2206 VSS.n1241 VSS.n1158 147.374
R2207 VSS.n1245 VSS.n1159 147.374
R2208 VSS.n1249 VSS.n1160 147.374
R2209 VSS.n1253 VSS.n1161 147.374
R2210 VSS.n1257 VSS.n1162 147.374
R2211 VSS.n1261 VSS.n1163 147.374
R2212 VSS.n1265 VSS.n1164 147.374
R2213 VSS.n1269 VSS.n1165 147.374
R2214 VSS.n1273 VSS.n1166 147.374
R2215 VSS.n1277 VSS.n1167 147.374
R2216 VSS.n1281 VSS.n1168 147.374
R2217 VSS.n1289 VSS.n1170 147.374
R2218 VSS.n1293 VSS.n1171 147.374
R2219 VSS.n1297 VSS.n1172 147.374
R2220 VSS.n1301 VSS.n1173 147.374
R2221 VSS.n1305 VSS.n1174 147.374
R2222 VSS.n1309 VSS.n1175 147.374
R2223 VSS.n1313 VSS.n1176 147.374
R2224 VSS.n1317 VSS.n1177 147.374
R2225 VSS.n1321 VSS.n1178 147.374
R2226 VSS.n1325 VSS.n1179 147.374
R2227 VSS.n1329 VSS.n1180 147.374
R2228 VSS.n1337 VSS.n1182 147.374
R2229 VSS.n1341 VSS.n1183 147.374
R2230 VSS.n1345 VSS.n1184 147.374
R2231 VSS.n1349 VSS.n1185 147.374
R2232 VSS.n1353 VSS.n1186 147.374
R2233 VSS.n1357 VSS.n1187 147.374
R2234 VSS.n1361 VSS.n1188 147.374
R2235 VSS.n1365 VSS.n1189 147.374
R2236 VSS.n1191 VSS.n1190 147.374
R2237 VSS.n1371 VSS.n1155 147.374
R2238 VSS.n1373 VSS.n1152 147.374
R2239 VSS.n2014 VSS.n788 147.374
R2240 VSS.n2009 VSS.n790 147.374
R2241 VSS.n2006 VSS.n791 147.374
R2242 VSS.n2002 VSS.n792 147.374
R2243 VSS.n1998 VSS.n793 147.374
R2244 VSS.n1994 VSS.n794 147.374
R2245 VSS.n1990 VSS.n795 147.374
R2246 VSS.n1986 VSS.n796 147.374
R2247 VSS.n1982 VSS.n797 147.374
R2248 VSS.n1976 VSS.n1975 147.374
R2249 VSS.n842 VSS.n803 147.374
R2250 VSS.n1968 VSS.n804 147.374
R2251 VSS.n1964 VSS.n805 147.374
R2252 VSS.n1960 VSS.n806 147.374
R2253 VSS.n1956 VSS.n807 147.374
R2254 VSS.n1952 VSS.n808 147.374
R2255 VSS.n1948 VSS.n809 147.374
R2256 VSS.n1944 VSS.n810 147.374
R2257 VSS.n1940 VSS.n811 147.374
R2258 VSS.n1936 VSS.n812 147.374
R2259 VSS.n1932 VSS.n813 147.374
R2260 VSS.n1928 VSS.n814 147.374
R2261 VSS.n1924 VSS.n815 147.374
R2262 VSS.n1920 VSS.n816 147.374
R2263 VSS.n1916 VSS.n817 147.374
R2264 VSS.n1912 VSS.n818 147.374
R2265 VSS.n1908 VSS.n819 147.374
R2266 VSS.n1904 VSS.n820 147.374
R2267 VSS.n1900 VSS.n821 147.374
R2268 VSS.n1896 VSS.n822 147.374
R2269 VSS.n1892 VSS.n823 147.374
R2270 VSS.n1888 VSS.n824 147.374
R2271 VSS.n1884 VSS.n825 147.374
R2272 VSS.n1880 VSS.n826 147.374
R2273 VSS.n1876 VSS.n827 147.374
R2274 VSS.n1872 VSS.n828 147.374
R2275 VSS.n1868 VSS.n829 147.374
R2276 VSS.n1864 VSS.n830 147.374
R2277 VSS.n1860 VSS.n831 147.374
R2278 VSS.n1856 VSS.n832 147.374
R2279 VSS.n1852 VSS.n833 147.374
R2280 VSS.n1848 VSS.n834 147.374
R2281 VSS.n1844 VSS.n835 147.374
R2282 VSS.n1840 VSS.n836 147.374
R2283 VSS.n1836 VSS.n837 147.374
R2284 VSS.n545 VSS.n544 147.374
R2285 VSS.n546 VSS.n540 147.374
R2286 VSS.n2097 VSS.n2096 147.374
R2287 VSS.n635 VSS.n522 147.374
R2288 VSS.n547 VSS.n546 147.374
R2289 VSS.n544 VSS.n543 147.374
R2290 VSS.n2098 VSS.n2097 147.374
R2291 VSS.n635 VSS.n634 147.374
R2292 VSS.n2014 VSS.n2013 147.374
R2293 VSS.n2007 VSS.n790 147.374
R2294 VSS.n2003 VSS.n791 147.374
R2295 VSS.n1999 VSS.n792 147.374
R2296 VSS.n1995 VSS.n793 147.374
R2297 VSS.n1991 VSS.n794 147.374
R2298 VSS.n1987 VSS.n795 147.374
R2299 VSS.n1983 VSS.n796 147.374
R2300 VSS.n1979 VSS.n797 147.374
R2301 VSS.n1226 VSS.n645 147.374
R2302 VSS.n1222 VSS.n644 147.374
R2303 VSS.n1218 VSS.n643 147.374
R2304 VSS.n1214 VSS.n642 147.374
R2305 VSS.n1210 VSS.n641 147.374
R2306 VSS.n1206 VSS.n640 147.374
R2307 VSS.n1202 VSS.n639 147.374
R2308 VSS.n1198 VSS.n638 147.374
R2309 VSS.n1194 VSS.n637 147.374
R2310 VSS.n647 VSS.n636 147.374
R2311 VSS.n1539 VSS.n1118 147.374
R2312 VSS.n1531 VSS.n1107 147.374
R2313 VSS.n1527 VSS.n1108 147.374
R2314 VSS.n1523 VSS.n1109 147.374
R2315 VSS.n1519 VSS.n1110 147.374
R2316 VSS.n1515 VSS.n1111 147.374
R2317 VSS.n1511 VSS.n1112 147.374
R2318 VSS.n1507 VSS.n1113 147.374
R2319 VSS.n1503 VSS.n1114 147.374
R2320 VSS.n1499 VSS.n1115 147.374
R2321 VSS.n1495 VSS.n1116 147.374
R2322 VSS.n1413 VSS.n1412 147.374
R2323 VSS.n1409 VSS.n1407 147.374
R2324 VSS.n1420 VSS.n1419 147.374
R2325 VSS.n1406 VSS.n1404 147.374
R2326 VSS.n1427 VSS.n1426 147.374
R2327 VSS.n1403 VSS.n1401 147.374
R2328 VSS.n1434 VSS.n1433 147.374
R2329 VSS.n1400 VSS.n1398 147.374
R2330 VSS.n1441 VSS.n1440 147.374
R2331 VSS.n1397 VSS.n1395 147.374
R2332 VSS.n1448 VSS.n1447 147.374
R2333 VSS.n1813 VSS.n1812 147.374
R2334 VSS.n1807 VSS.n859 147.374
R2335 VSS.n1805 VSS.n1804 147.374
R2336 VSS.n1800 VSS.n1799 147.374
R2337 VSS.n1797 VSS.n1796 147.374
R2338 VSS.n1790 VSS.n1789 147.374
R2339 VSS.n1787 VSS.n1786 147.374
R2340 VSS.n1782 VSS.n1781 147.374
R2341 VSS.n1779 VSS.n1778 147.374
R2342 VSS.n1774 VSS.n1773 147.374
R2343 VSS.n1771 VSS.n1770 147.374
R2344 VSS.n1695 VSS.n1675 147.374
R2345 VSS.n1699 VSS.n1676 147.374
R2346 VSS.n1703 VSS.n1677 147.374
R2347 VSS.n1707 VSS.n1678 147.374
R2348 VSS.n1711 VSS.n1679 147.374
R2349 VSS.n1715 VSS.n1680 147.374
R2350 VSS.n1719 VSS.n1681 147.374
R2351 VSS.n1723 VSS.n1682 147.374
R2352 VSS.n1727 VSS.n1683 147.374
R2353 VSS.n1731 VSS.n1684 147.374
R2354 VSS.n1686 VSS.n1685 147.374
R2355 VSS.n2449 VSS.n100 147.374
R2356 VSS.n2441 VSS.n81 147.374
R2357 VSS.n2437 VSS.n82 147.374
R2358 VSS.n2433 VSS.n83 147.374
R2359 VSS.n2429 VSS.n84 147.374
R2360 VSS.n2425 VSS.n85 147.374
R2361 VSS.n2421 VSS.n86 147.374
R2362 VSS.n2417 VSS.n87 147.374
R2363 VSS.n2413 VSS.n88 147.374
R2364 VSS.n2402 VSS.n89 147.374
R2365 VSS.n2406 VSS.n90 147.374
R2366 VSS.n2452 VSS.n2451 147.374
R2367 VSS.n2369 VSS.n91 147.374
R2368 VSS.n2373 VSS.n92 147.374
R2369 VSS.n2377 VSS.n93 147.374
R2370 VSS.n2381 VSS.n94 147.374
R2371 VSS.n2385 VSS.n95 147.374
R2372 VSS.n2389 VSS.n96 147.374
R2373 VSS.n2392 VSS.n97 147.374
R2374 VSS.n418 VSS.n417 147.374
R2375 VSS.n415 VSS.n414 147.374
R2376 VSS.n410 VSS.n409 147.374
R2377 VSS.n407 VSS.n406 147.374
R2378 VSS.n402 VSS.n401 147.374
R2379 VSS.n399 VSS.n398 147.374
R2380 VSS.n394 VSS.n393 147.374
R2381 VSS.n391 VSS.n390 147.374
R2382 VSS.n283 VSS.n282 147.374
R2383 VSS.n280 VSS.n279 147.374
R2384 VSS.n275 VSS.n274 147.374
R2385 VSS.n272 VSS.n271 147.374
R2386 VSS.n267 VSS.n266 147.374
R2387 VSS.n264 VSS.n263 147.374
R2388 VSS.n259 VSS.n258 147.374
R2389 VSS.n256 VSS.n255 147.374
R2390 VSS.n251 VSS.n250 147.374
R2391 VSS.n248 VSS.n247 147.374
R2392 VSS.n243 VSS.n242 147.374
R2393 VSS.n1975 VSS.n801 147.374
R2394 VSS.n1969 VSS.n803 147.374
R2395 VSS.n1965 VSS.n804 147.374
R2396 VSS.n1961 VSS.n805 147.374
R2397 VSS.n1957 VSS.n806 147.374
R2398 VSS.n1953 VSS.n807 147.374
R2399 VSS.n1949 VSS.n808 147.374
R2400 VSS.n1945 VSS.n809 147.374
R2401 VSS.n1941 VSS.n810 147.374
R2402 VSS.n1937 VSS.n811 147.374
R2403 VSS.n1933 VSS.n812 147.374
R2404 VSS.n1929 VSS.n813 147.374
R2405 VSS.n1925 VSS.n814 147.374
R2406 VSS.n1921 VSS.n815 147.374
R2407 VSS.n1917 VSS.n816 147.374
R2408 VSS.n1913 VSS.n817 147.374
R2409 VSS.n1909 VSS.n818 147.374
R2410 VSS.n1905 VSS.n819 147.374
R2411 VSS.n1901 VSS.n820 147.374
R2412 VSS.n1897 VSS.n821 147.374
R2413 VSS.n1893 VSS.n822 147.374
R2414 VSS.n1889 VSS.n823 147.374
R2415 VSS.n1885 VSS.n824 147.374
R2416 VSS.n1881 VSS.n825 147.374
R2417 VSS.n1877 VSS.n826 147.374
R2418 VSS.n1873 VSS.n827 147.374
R2419 VSS.n1869 VSS.n828 147.374
R2420 VSS.n1865 VSS.n829 147.374
R2421 VSS.n1861 VSS.n830 147.374
R2422 VSS.n1857 VSS.n831 147.374
R2423 VSS.n1853 VSS.n832 147.374
R2424 VSS.n1849 VSS.n833 147.374
R2425 VSS.n1845 VSS.n834 147.374
R2426 VSS.n1841 VSS.n835 147.374
R2427 VSS.n1837 VSS.n836 147.374
R2428 VSS.n1833 VSS.n837 147.374
R2429 VSS.n1374 VSS.n1373 147.374
R2430 VSS.n1371 VSS.n1370 147.374
R2431 VSS.n1366 VSS.n1190 147.374
R2432 VSS.n1362 VSS.n1189 147.374
R2433 VSS.n1358 VSS.n1188 147.374
R2434 VSS.n1354 VSS.n1187 147.374
R2435 VSS.n1350 VSS.n1186 147.374
R2436 VSS.n1346 VSS.n1185 147.374
R2437 VSS.n1342 VSS.n1184 147.374
R2438 VSS.n1338 VSS.n1183 147.374
R2439 VSS.n1334 VSS.n1182 147.374
R2440 VSS.n1326 VSS.n1180 147.374
R2441 VSS.n1322 VSS.n1179 147.374
R2442 VSS.n1318 VSS.n1178 147.374
R2443 VSS.n1314 VSS.n1177 147.374
R2444 VSS.n1310 VSS.n1176 147.374
R2445 VSS.n1306 VSS.n1175 147.374
R2446 VSS.n1302 VSS.n1174 147.374
R2447 VSS.n1298 VSS.n1173 147.374
R2448 VSS.n1294 VSS.n1172 147.374
R2449 VSS.n1290 VSS.n1171 147.374
R2450 VSS.n1286 VSS.n1170 147.374
R2451 VSS.n1278 VSS.n1168 147.374
R2452 VSS.n1274 VSS.n1167 147.374
R2453 VSS.n1270 VSS.n1166 147.374
R2454 VSS.n1266 VSS.n1165 147.374
R2455 VSS.n1262 VSS.n1164 147.374
R2456 VSS.n1258 VSS.n1163 147.374
R2457 VSS.n1254 VSS.n1162 147.374
R2458 VSS.n1250 VSS.n1161 147.374
R2459 VSS.n1246 VSS.n1160 147.374
R2460 VSS.n1242 VSS.n1159 147.374
R2461 VSS.n1238 VSS.n1158 147.374
R2462 VSS.n1230 VSS.n1156 147.374
R2463 VSS.n1666 VSS.n1665 147.374
R2464 VSS.n1660 VSS.n889 147.374
R2465 VSS.n1657 VSS.n890 147.374
R2466 VSS.n1653 VSS.n891 147.374
R2467 VSS.n1649 VSS.n892 147.374
R2468 VSS.n1645 VSS.n893 147.374
R2469 VSS.n1641 VSS.n894 147.374
R2470 VSS.n1637 VSS.n895 147.374
R2471 VSS.n1633 VSS.n896 147.374
R2472 VSS.n1629 VSS.n897 147.374
R2473 VSS.n1625 VSS.n898 147.374
R2474 VSS.n1551 VSS.n1049 147.374
R2475 VSS.n1054 VSS.n1053 147.374
R2476 VSS.n1066 VSS.n1055 147.374
R2477 VSS.n1070 VSS.n1056 147.374
R2478 VSS.n1074 VSS.n1057 147.374
R2479 VSS.n1078 VSS.n1058 147.374
R2480 VSS.n1082 VSS.n1059 147.374
R2481 VSS.n1086 VSS.n1060 147.374
R2482 VSS.n1090 VSS.n1061 147.374
R2483 VSS.n1094 VSS.n1062 147.374
R2484 VSS.n1101 VSS.n1063 147.374
R2485 VSS.n1101 VSS.n1100 147.374
R2486 VSS.n1096 VSS.n1062 147.374
R2487 VSS.n1093 VSS.n1061 147.374
R2488 VSS.n1089 VSS.n1060 147.374
R2489 VSS.n1085 VSS.n1059 147.374
R2490 VSS.n1081 VSS.n1058 147.374
R2491 VSS.n1077 VSS.n1057 147.374
R2492 VSS.n1073 VSS.n1056 147.374
R2493 VSS.n1069 VSS.n1055 147.374
R2494 VSS.n1065 VSS.n1054 147.374
R2495 VSS.n1552 VSS.n1551 147.374
R2496 VSS.n1666 VSS.n900 147.374
R2497 VSS.n1658 VSS.n889 147.374
R2498 VSS.n1654 VSS.n890 147.374
R2499 VSS.n1650 VSS.n891 147.374
R2500 VSS.n1646 VSS.n892 147.374
R2501 VSS.n1642 VSS.n893 147.374
R2502 VSS.n1638 VSS.n894 147.374
R2503 VSS.n1634 VSS.n895 147.374
R2504 VSS.n1630 VSS.n896 147.374
R2505 VSS.n1626 VSS.n897 147.374
R2506 VSS.n1622 VSS.n898 147.374
R2507 VSS.n70 VSS.n46 140.69
R2508 VSS.n63 VSS.n46 140.69
R2509 VSS.n17 VSS.n16 140.69
R2510 VSS.n17 VSS.n8 140.69
R2511 VSS.n750 VSS.n749 140.69
R2512 VSS.n749 VSS.n723 140.69
R2513 VSS.n742 VSS.n723 140.69
R2514 VSS.n742 VSS.n741 140.69
R2515 VSS.n741 VSS.n727 140.69
R2516 VSS.n734 VSS.n727 140.69
R2517 VSS.n734 VSS.n733 140.69
R2518 VSS.n690 VSS.n684 140.69
R2519 VSS.n697 VSS.n684 140.69
R2520 VSS.n698 VSS.n697 140.69
R2521 VSS.n698 VSS.n680 140.69
R2522 VSS.n706 VSS.n680 140.69
R2523 VSS.n707 VSS.n706 140.69
R2524 VSS.n707 VSS.n677 140.69
R2525 VSS.n999 VSS.n993 140.69
R2526 VSS.n1000 VSS.n999 140.69
R2527 VSS.n1000 VSS.n989 140.69
R2528 VSS.n1007 VSS.n989 140.69
R2529 VSS.n1008 VSS.n1007 140.69
R2530 VSS.n1008 VSS.n985 140.69
R2531 VSS.n1015 VSS.n985 140.69
R2532 VSS.n974 VSS.n941 140.69
R2533 VSS.n967 VSS.n941 140.69
R2534 VSS.n967 VSS.n966 140.69
R2535 VSS.n966 VSS.n945 140.69
R2536 VSS.n959 VSS.n945 140.69
R2537 VSS.n959 VSS.n958 140.69
R2538 VSS.n958 VSS.n949 140.69
R2539 VSS.n2156 VSS.n2155 117.233
R2540 VSS.n552 VSS.n535 99.5348
R2541 VSS.n558 VSS.n535 99.5348
R2542 VSS.n558 VSS.n531 99.5348
R2543 VSS.n565 VSS.n531 99.5348
R2544 VSS.n565 VSS.n527 99.5348
R2545 VSS.n571 VSS.n527 99.5348
R2546 VSS.n571 VSS.n435 99.5348
R2547 VSS.n2195 VSS.n437 99.5348
R2548 VSS.n2189 VSS.n437 99.5348
R2549 VSS.n2189 VSS.n2188 99.5348
R2550 VSS.n2188 VSS.n2187 99.5348
R2551 VSS.n2187 VSS.n446 99.5348
R2552 VSS.n2181 VSS.n446 99.5348
R2553 VSS.n2181 VSS.n2180 99.5348
R2554 VSS.n2180 VSS.n2179 99.5348
R2555 VSS.n2179 VSS.n453 99.5348
R2556 VSS.n2173 VSS.n453 99.5348
R2557 VSS.n2173 VSS.n2172 99.5348
R2558 VSS.n2172 VSS.n2171 99.5348
R2559 VSS.n2171 VSS.n460 99.5348
R2560 VSS.n2165 VSS.n460 99.5348
R2561 VSS.n2165 VSS.n2164 99.5348
R2562 VSS.n2164 VSS.n2163 99.5348
R2563 VSS.n2163 VSS.n467 99.5348
R2564 VSS.n2157 VSS.n467 99.5348
R2565 VSS.n2093 VSS.n646 99.5348
R2566 VSS.n2087 VSS.n2086 99.5348
R2567 VSS.n2086 VSS.n2085 99.5348
R2568 VSS.n2085 VSS.n652 99.5348
R2569 VSS.n2079 VSS.n2078 99.5348
R2570 VSS.n2078 VSS.n2077 99.5348
R2571 VSS.n2077 VSS.n656 99.5348
R2572 VSS.n2071 VSS.n2070 99.5348
R2573 VSS.n2070 VSS.n2069 99.5348
R2574 VSS.n2069 VSS.n660 99.5348
R2575 VSS.n2063 VSS.n2062 99.5348
R2576 VSS.n2062 VSS.n2061 99.5348
R2577 VSS.n1043 VSS.n1036 99.5348
R2578 VSS.n1037 VSS.n1036 99.5348
R2579 VSS.n2048 VSS.n772 99.5348
R2580 VSS.n2048 VSS.n2047 99.5348
R2581 VSS.n2047 VSS.n2046 99.5348
R2582 VSS.n2040 VSS.n777 99.5348
R2583 VSS.n2040 VSS.n2039 99.5348
R2584 VSS.n2039 VSS.n2038 99.5348
R2585 VSS.n2032 VSS.n781 99.5348
R2586 VSS.n2032 VSS.n2031 99.5348
R2587 VSS.n2031 VSS.n2030 99.5348
R2588 VSS.n2024 VSS.n785 99.5348
R2589 VSS.n2024 VSS.n2023 99.5348
R2590 VSS.n2023 VSS.n2022 99.5348
R2591 VSS.n2016 VSS.n789 99.5348
R2592 VSS.t36 VSS.n646 92.2161
R2593 VSS.n789 VSS.t19 92.2161
R2594 VSS.n313 VSS.t57 90.6265
R2595 VSS.n297 VSS.t49 90.6265
R2596 VSS.n369 VSS.t67 90.6265
R2597 VSS.n352 VSS.t60 90.6265
R2598 VSS.t79 VSS.n1043 89.2886
R2599 VSS.n1037 VSS.t13 89.2886
R2600 VSS.n554 VSS.n537 85.8358
R2601 VSS.n550 VSS.n549 85.8358
R2602 VSS.n633 VSS.n632 85.8358
R2603 VSS.n1451 VSS.n1450 82.4476
R2604 VSS.n1537 VSS.n1120 82.4476
R2605 VSS.n1410 VSS.n1148 82.4476
R2606 VSS.n1496 VSS.n1121 82.4476
R2607 VSS.n1735 VSS.n875 82.4476
R2608 VSS.n1816 VSS.n1815 82.4476
R2609 VSS.n1693 VSS.n1689 82.4476
R2610 VSS.n1769 VSS.n1768 82.4476
R2611 VSS.n1556 VSS.n1554 82.4476
R2612 VSS.n1560 VSS.n1045 82.4476
R2613 VSS.n1664 VSS.n902 82.4476
R2614 VSS.n1623 VSS.n903 82.4476
R2615 VSS.n313 VSS.t55 81.8918
R2616 VSS.n312 VSS.t99 81.8918
R2617 VSS.n297 VSS.t46 81.8918
R2618 VSS.n373 VSS.t64 81.8918
R2619 VSS.n369 VSS.t66 81.8918
R2620 VSS.n352 VSS.t58 81.8918
R2621 VSS.n48 VSS.t61 81.8918
R2622 VSS.n61 VSS.t86 81.8918
R2623 VSS.n7 VSS.t97 81.8918
R2624 VSS.n24 VSS.t95 81.8918
R2625 VSS.n2061 VSS.n664 79.0424
R2626 VSS.n425 VSS.n218 76.8005
R2627 VSS.n2447 VSS.n2400 76.8005
R2628 VSS.n421 VSS.n420 76.8005
R2629 VSS.n2394 VSS.n2393 76.8005
R2630 VSS.n2018 VSS.n787 76.8005
R2631 VSS.n1832 VSS.n1831 76.8005
R2632 VSS.n1390 VSS.n1376 76.8005
R2633 VSS.n2091 VSS.n649 76.8005
R2634 VSS.n2197 VSS.n435 74.6512
R2635 VSS.t39 VSS.n652 71.7237
R2636 VSS.n785 VSS.t12 71.7237
R2637 VSS.n63 VSS.t88 70.3453
R2638 VSS.t98 VSS.n8 70.3453
R2639 VSS.n733 VSS.t83 70.3453
R2640 VSS.t37 VSS.n677 70.3453
R2641 VSS.t43 VSS.n993 70.3453
R2642 VSS.t45 VSS.n974 70.3453
R2643 VSS.n2063 VSS.t9 68.7962
R2644 VSS.n2046 VSS.t51 68.7962
R2645 VSS.n1818 VSS.n855 66.162
R2646 VSS.n1972 VSS.n1971 64.7534
R2647 VSS.n1236 VSS.n1235 64.7534
R2648 VSS.n2104 VSS.n2103 62.1181
R2649 VSS.n1372 VSS.n98 61.9943
R2650 VSS.n423 VSS.n220 54.18
R2651 VSS.n2450 VSS.n80 54.18
R2652 VSS.t10 VSS.n656 51.2314
R2653 VSS.n781 VSS.t2 51.2314
R2654 VSS.n2157 VSS.t128 49.7676
R2655 VSS.n2071 VSS.t10 48.3039
R2656 VSS.n2038 VSS.t2 48.3039
R2657 VSS.n1926 VSS.n1923 39.1534
R2658 VSS.n1878 VSS.n1875 39.1534
R2659 VSS.n1284 VSS.n1283 39.1534
R2660 VSS.n1332 VSS.n1331 39.1534
R2661 VSS.t128 VSS.n2156 38.2032
R2662 VSS.n423 VSS.n216 35.4256
R2663 VSS.n429 VSS.n216 35.4256
R2664 VSS.n2198 VSS.n212 35.4256
R2665 VSS.n2204 VSS.n205 35.4256
R2666 VSS.n2211 VSS.n205 35.4256
R2667 VSS.n2211 VSS.n2210 35.4256
R2668 VSS.n2217 VSS.n198 35.4256
R2669 VSS.n2224 VSS.n198 35.4256
R2670 VSS.n2224 VSS.n2223 35.4256
R2671 VSS.n2230 VSS.n191 35.4256
R2672 VSS.n2237 VSS.n191 35.4256
R2673 VSS.n2237 VSS.n2236 35.4256
R2674 VSS.n2243 VSS.n184 35.4256
R2675 VSS.n2250 VSS.n184 35.4256
R2676 VSS.n2250 VSS.n2249 35.4256
R2677 VSS.n2256 VSS.n177 35.4256
R2678 VSS.n2262 VSS.n177 35.4256
R2679 VSS.n2268 VSS.n173 35.4256
R2680 VSS.n2268 VSS.n169 35.4256
R2681 VSS.n2274 VSS.n169 35.4256
R2682 VSS.n2280 VSS.n165 35.4256
R2683 VSS.n2280 VSS.n161 35.4256
R2684 VSS.n2286 VSS.n161 35.4256
R2685 VSS.n2292 VSS.n157 35.4256
R2686 VSS.n2292 VSS.n153 35.4256
R2687 VSS.n2298 VSS.n153 35.4256
R2688 VSS.n2304 VSS.n148 35.4256
R2689 VSS.n2304 VSS.n149 35.4256
R2690 VSS.n2310 VSS.n140 35.4256
R2691 VSS.n2316 VSS.n140 35.4256
R2692 VSS.n2316 VSS.n141 35.4256
R2693 VSS.n2322 VSS.n132 35.4256
R2694 VSS.n2328 VSS.n132 35.4256
R2695 VSS.n2328 VSS.n133 35.4256
R2696 VSS.n2334 VSS.n124 35.4256
R2697 VSS.n2340 VSS.n124 35.4256
R2698 VSS.n2340 VSS.n125 35.4256
R2699 VSS.n2346 VSS.n116 35.4256
R2700 VSS.n2352 VSS.n116 35.4256
R2701 VSS.n2352 VSS.n117 35.4256
R2702 VSS.n2358 VSS.n109 35.4256
R2703 VSS.n2364 VSS.n109 35.4256
R2704 VSS.n2397 VSS.n104 35.4256
R2705 VSS.n2397 VSS.n80 35.4256
R2706 VSS.n1454 VSS.n1150 35.4256
R2707 VSS.n1125 VSS.n1106 35.4256
R2708 VSS.n1542 VSS.n1541 35.4256
R2709 VSS.n1549 VSS.n1047 35.4256
R2710 VSS.n1668 VSS.n888 35.4256
R2711 VSS.n1674 VSS.n884 35.4256
R2712 VSS.n1739 VSS.n1738 35.4256
R2713 VSS.n1974 VSS.n802 35.4256
R2714 VSS.n1974 VSS.n840 35.4256
R2715 VSS.n1820 VSS.n840 35.4256
R2716 VSS.n1819 VSS.n1818 35.4256
R2717 VSS.n2256 VSS.t28 34.9046
R2718 VSS.n149 VSS.t15 34.9046
R2719 VSS.t59 VSS.n212 33.8627
R2720 VSS.n2364 VSS.t47 33.8627
R2721 VSS.n304 VSS.n303 32.8962
R2722 VSS.n359 VSS.n358 32.8962
R2723 VSS.t9 VSS.n660 30.739
R2724 VSS.n777 VSS.t51 30.739
R2725 VSS.n2197 VSS.n2196 30.7369
R2726 VSS.n2196 VSS.t20 29.695
R2727 VSS.n2358 VSS.t62 29.695
R2728 VSS.n2262 VSS.t5 28.6531
R2729 VSS.t31 VSS.n148 28.6531
R2730 VSS.n64 VSS.n62 28.3989
R2731 VSS.n21 VSS.n20 28.3989
R2732 VSS.n328 VSS.n327 27.9576
R2733 VSS.n332 VSS.n331 27.9576
R2734 VSS.n336 VSS.n335 27.9576
R2735 VSS.n340 VSS.n339 27.9576
R2736 VSS.n344 VSS.n343 27.9576
R2737 VSS.n2079 VSS.t39 27.8115
R2738 VSS.n2030 VSS.t12 27.8115
R2739 VSS.n326 VSS.n325 27.7293
R2740 VSS.n330 VSS.n329 27.7293
R2741 VSS.n334 VSS.n333 27.7293
R2742 VSS.n338 VSS.n337 27.7293
R2743 VSS.n342 VSS.n341 27.7293
R2744 VSS.n346 VSS.n345 27.7293
R2745 VSS.n42 VSS.n41 27.7293
R2746 VSS.n40 VSS.n39 27.7293
R2747 VSS.n38 VSS.n37 27.7293
R2748 VSS.n36 VSS.n35 27.7293
R2749 VSS.n34 VSS.n33 27.7293
R2750 VSS.n2243 VSS.t25 27.6112
R2751 VSS.n141 VSS.t3 27.6112
R2752 VSS.n1737 VSS.n1674 27.6112
R2753 VSS.n320 VSS.n291 27.5286
R2754 VSS.n321 VSS.n289 27.5286
R2755 VSS.n381 VSS.n364 27.5286
R2756 VSS.n380 VSS.n366 27.5286
R2757 VSS.n58 VSS.n49 27.5286
R2758 VSS.n29 VSS.n6 27.5286
R2759 VSS.n754 VSS.n720 25.6009
R2760 VSS.n689 VSS.n688 25.6009
R2761 VSS.n1017 VSS.n1016 25.6009
R2762 VSS.n952 VSS.n951 25.6009
R2763 VSS.n426 VSS.n425 25.6005
R2764 VSS.n427 VSS.n426 25.6005
R2765 VSS.n427 VSS.n210 25.6005
R2766 VSS.n2200 VSS.n210 25.6005
R2767 VSS.n2201 VSS.n2200 25.6005
R2768 VSS.n2202 VSS.n2201 25.6005
R2769 VSS.n2202 VSS.n203 25.6005
R2770 VSS.n2213 VSS.n203 25.6005
R2771 VSS.n2214 VSS.n2213 25.6005
R2772 VSS.n2215 VSS.n2214 25.6005
R2773 VSS.n2215 VSS.n196 25.6005
R2774 VSS.n2226 VSS.n196 25.6005
R2775 VSS.n2227 VSS.n2226 25.6005
R2776 VSS.n2228 VSS.n2227 25.6005
R2777 VSS.n2228 VSS.n189 25.6005
R2778 VSS.n2239 VSS.n189 25.6005
R2779 VSS.n2240 VSS.n2239 25.6005
R2780 VSS.n2241 VSS.n2240 25.6005
R2781 VSS.n2241 VSS.n182 25.6005
R2782 VSS.n2252 VSS.n182 25.6005
R2783 VSS.n2253 VSS.n2252 25.6005
R2784 VSS.n2254 VSS.n2253 25.6005
R2785 VSS.n2254 VSS.n175 25.6005
R2786 VSS.n2264 VSS.n175 25.6005
R2787 VSS.n2265 VSS.n2264 25.6005
R2788 VSS.n2266 VSS.n2265 25.6005
R2789 VSS.n2266 VSS.n167 25.6005
R2790 VSS.n2276 VSS.n167 25.6005
R2791 VSS.n2277 VSS.n2276 25.6005
R2792 VSS.n2278 VSS.n2277 25.6005
R2793 VSS.n2278 VSS.n159 25.6005
R2794 VSS.n2288 VSS.n159 25.6005
R2795 VSS.n2289 VSS.n2288 25.6005
R2796 VSS.n2290 VSS.n2289 25.6005
R2797 VSS.n2290 VSS.n151 25.6005
R2798 VSS.n2300 VSS.n151 25.6005
R2799 VSS.n2301 VSS.n2300 25.6005
R2800 VSS.n2302 VSS.n2301 25.6005
R2801 VSS.n2302 VSS.n143 25.6005
R2802 VSS.n2312 VSS.n143 25.6005
R2803 VSS.n2313 VSS.n2312 25.6005
R2804 VSS.n2314 VSS.n2313 25.6005
R2805 VSS.n2314 VSS.n135 25.6005
R2806 VSS.n2324 VSS.n135 25.6005
R2807 VSS.n2325 VSS.n2324 25.6005
R2808 VSS.n2326 VSS.n2325 25.6005
R2809 VSS.n2326 VSS.n127 25.6005
R2810 VSS.n2336 VSS.n127 25.6005
R2811 VSS.n2337 VSS.n2336 25.6005
R2812 VSS.n2338 VSS.n2337 25.6005
R2813 VSS.n2338 VSS.n119 25.6005
R2814 VSS.n2348 VSS.n119 25.6005
R2815 VSS.n2349 VSS.n2348 25.6005
R2816 VSS.n2350 VSS.n2349 25.6005
R2817 VSS.n2350 VSS.n111 25.6005
R2818 VSS.n2360 VSS.n111 25.6005
R2819 VSS.n2361 VSS.n2360 25.6005
R2820 VSS.n2362 VSS.n2361 25.6005
R2821 VSS.n2362 VSS.n102 25.6005
R2822 VSS.n2399 VSS.n102 25.6005
R2823 VSS.n2400 VSS.n2399 25.6005
R2824 VSS.n244 VSS.n218 25.6005
R2825 VSS.n245 VSS.n244 25.6005
R2826 VSS.n246 VSS.n245 25.6005
R2827 VSS.n246 VSS.n240 25.6005
R2828 VSS.n252 VSS.n240 25.6005
R2829 VSS.n253 VSS.n252 25.6005
R2830 VSS.n254 VSS.n253 25.6005
R2831 VSS.n254 VSS.n238 25.6005
R2832 VSS.n260 VSS.n238 25.6005
R2833 VSS.n261 VSS.n260 25.6005
R2834 VSS.n262 VSS.n261 25.6005
R2835 VSS.n262 VSS.n236 25.6005
R2836 VSS.n268 VSS.n236 25.6005
R2837 VSS.n269 VSS.n268 25.6005
R2838 VSS.n270 VSS.n269 25.6005
R2839 VSS.n270 VSS.n234 25.6005
R2840 VSS.n276 VSS.n234 25.6005
R2841 VSS.n277 VSS.n276 25.6005
R2842 VSS.n278 VSS.n277 25.6005
R2843 VSS.n284 VSS.n232 25.6005
R2844 VSS.n389 VSS.n228 25.6005
R2845 VSS.n395 VSS.n228 25.6005
R2846 VSS.n396 VSS.n395 25.6005
R2847 VSS.n397 VSS.n396 25.6005
R2848 VSS.n397 VSS.n226 25.6005
R2849 VSS.n403 VSS.n226 25.6005
R2850 VSS.n404 VSS.n403 25.6005
R2851 VSS.n405 VSS.n404 25.6005
R2852 VSS.n405 VSS.n224 25.6005
R2853 VSS.n411 VSS.n224 25.6005
R2854 VSS.n412 VSS.n411 25.6005
R2855 VSS.n413 VSS.n412 25.6005
R2856 VSS.n413 VSS.n222 25.6005
R2857 VSS.n419 VSS.n222 25.6005
R2858 VSS.n420 VSS.n419 25.6005
R2859 VSS.n421 VSS.n214 25.6005
R2860 VSS.n431 VSS.n214 25.6005
R2861 VSS.n432 VSS.n431 25.6005
R2862 VSS.n433 VSS.n432 25.6005
R2863 VSS.n433 VSS.n207 25.6005
R2864 VSS.n2206 VSS.n207 25.6005
R2865 VSS.n2207 VSS.n2206 25.6005
R2866 VSS.n2208 VSS.n2207 25.6005
R2867 VSS.n2208 VSS.n200 25.6005
R2868 VSS.n2219 VSS.n200 25.6005
R2869 VSS.n2220 VSS.n2219 25.6005
R2870 VSS.n2221 VSS.n2220 25.6005
R2871 VSS.n2221 VSS.n193 25.6005
R2872 VSS.n2232 VSS.n193 25.6005
R2873 VSS.n2233 VSS.n2232 25.6005
R2874 VSS.n2234 VSS.n2233 25.6005
R2875 VSS.n2234 VSS.n186 25.6005
R2876 VSS.n2245 VSS.n186 25.6005
R2877 VSS.n2246 VSS.n2245 25.6005
R2878 VSS.n2247 VSS.n2246 25.6005
R2879 VSS.n2247 VSS.n179 25.6005
R2880 VSS.n2258 VSS.n179 25.6005
R2881 VSS.n2259 VSS.n2258 25.6005
R2882 VSS.n2260 VSS.n2259 25.6005
R2883 VSS.n2260 VSS.n171 25.6005
R2884 VSS.n2270 VSS.n171 25.6005
R2885 VSS.n2271 VSS.n2270 25.6005
R2886 VSS.n2272 VSS.n2271 25.6005
R2887 VSS.n2272 VSS.n163 25.6005
R2888 VSS.n2282 VSS.n163 25.6005
R2889 VSS.n2283 VSS.n2282 25.6005
R2890 VSS.n2284 VSS.n2283 25.6005
R2891 VSS.n2284 VSS.n155 25.6005
R2892 VSS.n2294 VSS.n155 25.6005
R2893 VSS.n2295 VSS.n2294 25.6005
R2894 VSS.n2296 VSS.n2295 25.6005
R2895 VSS.n2296 VSS.n146 25.6005
R2896 VSS.n2306 VSS.n146 25.6005
R2897 VSS.n2307 VSS.n2306 25.6005
R2898 VSS.n2308 VSS.n2307 25.6005
R2899 VSS.n2308 VSS.n138 25.6005
R2900 VSS.n2318 VSS.n138 25.6005
R2901 VSS.n2319 VSS.n2318 25.6005
R2902 VSS.n2320 VSS.n2319 25.6005
R2903 VSS.n2320 VSS.n130 25.6005
R2904 VSS.n2330 VSS.n130 25.6005
R2905 VSS.n2331 VSS.n2330 25.6005
R2906 VSS.n2332 VSS.n2331 25.6005
R2907 VSS.n2332 VSS.n122 25.6005
R2908 VSS.n2342 VSS.n122 25.6005
R2909 VSS.n2343 VSS.n2342 25.6005
R2910 VSS.n2344 VSS.n2343 25.6005
R2911 VSS.n2344 VSS.n114 25.6005
R2912 VSS.n2354 VSS.n114 25.6005
R2913 VSS.n2355 VSS.n2354 25.6005
R2914 VSS.n2356 VSS.n2355 25.6005
R2915 VSS.n2356 VSS.n107 25.6005
R2916 VSS.n2366 VSS.n107 25.6005
R2917 VSS.n2367 VSS.n2366 25.6005
R2918 VSS.n2395 VSS.n2367 25.6005
R2919 VSS.n2395 VSS.n2394 25.6005
R2920 VSS.n2447 VSS.n2446 25.6005
R2921 VSS.n2446 VSS.n2445 25.6005
R2922 VSS.n2445 VSS.n2444 25.6005
R2923 VSS.n2444 VSS.n2442 25.6005
R2924 VSS.n2442 VSS.n2439 25.6005
R2925 VSS.n2439 VSS.n2438 25.6005
R2926 VSS.n2438 VSS.n2435 25.6005
R2927 VSS.n2435 VSS.n2434 25.6005
R2928 VSS.n2434 VSS.n2431 25.6005
R2929 VSS.n2431 VSS.n2430 25.6005
R2930 VSS.n2430 VSS.n2427 25.6005
R2931 VSS.n2427 VSS.n2426 25.6005
R2932 VSS.n2426 VSS.n2423 25.6005
R2933 VSS.n2423 VSS.n2422 25.6005
R2934 VSS.n2422 VSS.n2419 25.6005
R2935 VSS.n2419 VSS.n2418 25.6005
R2936 VSS.n2418 VSS.n2415 25.6005
R2937 VSS.n2415 VSS.n2414 25.6005
R2938 VSS.n2414 VSS.n2411 25.6005
R2939 VSS.n2404 VSS.n2401 25.6005
R2940 VSS.n2453 VSS.n76 25.6005
R2941 VSS.n2453 VSS.n77 25.6005
R2942 VSS.n2368 VSS.n77 25.6005
R2943 VSS.n2371 VSS.n2368 25.6005
R2944 VSS.n2372 VSS.n2371 25.6005
R2945 VSS.n2375 VSS.n2372 25.6005
R2946 VSS.n2376 VSS.n2375 25.6005
R2947 VSS.n2379 VSS.n2376 25.6005
R2948 VSS.n2380 VSS.n2379 25.6005
R2949 VSS.n2383 VSS.n2380 25.6005
R2950 VSS.n2384 VSS.n2383 25.6005
R2951 VSS.n2387 VSS.n2384 25.6005
R2952 VSS.n2388 VSS.n2387 25.6005
R2953 VSS.n2391 VSS.n2388 25.6005
R2954 VSS.n2393 VSS.n2391 25.6005
R2955 VSS.n1452 VSS.n1451 25.6005
R2956 VSS.n1452 VSS.n1144 25.6005
R2957 VSS.n1462 VSS.n1144 25.6005
R2958 VSS.n1463 VSS.n1462 25.6005
R2959 VSS.n1464 VSS.n1463 25.6005
R2960 VSS.n1464 VSS.n1135 25.6005
R2961 VSS.n1479 VSS.n1135 25.6005
R2962 VSS.n1480 VSS.n1479 25.6005
R2963 VSS.n1482 VSS.n1480 25.6005
R2964 VSS.n1482 VSS.n1481 25.6005
R2965 VSS.n1481 VSS.n1120 25.6005
R2966 VSS.n1450 VSS.n1394 25.6005
R2967 VSS.n1445 VSS.n1394 25.6005
R2968 VSS.n1445 VSS.n1444 25.6005
R2969 VSS.n1444 VSS.n1443 25.6005
R2970 VSS.n1443 VSS.n1396 25.6005
R2971 VSS.n1438 VSS.n1396 25.6005
R2972 VSS.n1438 VSS.n1437 25.6005
R2973 VSS.n1437 VSS.n1436 25.6005
R2974 VSS.n1436 VSS.n1399 25.6005
R2975 VSS.n1431 VSS.n1399 25.6005
R2976 VSS.n1431 VSS.n1430 25.6005
R2977 VSS.n1430 VSS.n1429 25.6005
R2978 VSS.n1429 VSS.n1402 25.6005
R2979 VSS.n1424 VSS.n1402 25.6005
R2980 VSS.n1424 VSS.n1423 25.6005
R2981 VSS.n1423 VSS.n1422 25.6005
R2982 VSS.n1422 VSS.n1405 25.6005
R2983 VSS.n1417 VSS.n1405 25.6005
R2984 VSS.n1417 VSS.n1416 25.6005
R2985 VSS.n1416 VSS.n1415 25.6005
R2986 VSS.n1415 VSS.n1408 25.6005
R2987 VSS.n1410 VSS.n1408 25.6005
R2988 VSS.n1456 VSS.n1148 25.6005
R2989 VSS.n1457 VSS.n1456 25.6005
R2990 VSS.n1458 VSS.n1457 25.6005
R2991 VSS.n1458 VSS.n1140 25.6005
R2992 VSS.n1468 VSS.n1140 25.6005
R2993 VSS.n1469 VSS.n1468 25.6005
R2994 VSS.n1475 VSS.n1469 25.6005
R2995 VSS.n1475 VSS.n1474 25.6005
R2996 VSS.n1472 VSS.n1471 25.6005
R2997 VSS.n1537 VSS.n1536 25.6005
R2998 VSS.n1536 VSS.n1535 25.6005
R2999 VSS.n1535 VSS.n1534 25.6005
R3000 VSS.n1534 VSS.n1532 25.6005
R3001 VSS.n1532 VSS.n1529 25.6005
R3002 VSS.n1529 VSS.n1528 25.6005
R3003 VSS.n1528 VSS.n1525 25.6005
R3004 VSS.n1525 VSS.n1524 25.6005
R3005 VSS.n1524 VSS.n1521 25.6005
R3006 VSS.n1521 VSS.n1520 25.6005
R3007 VSS.n1520 VSS.n1517 25.6005
R3008 VSS.n1517 VSS.n1516 25.6005
R3009 VSS.n1516 VSS.n1513 25.6005
R3010 VSS.n1513 VSS.n1512 25.6005
R3011 VSS.n1512 VSS.n1509 25.6005
R3012 VSS.n1509 VSS.n1508 25.6005
R3013 VSS.n1508 VSS.n1505 25.6005
R3014 VSS.n1505 VSS.n1504 25.6005
R3015 VSS.n1504 VSS.n1501 25.6005
R3016 VSS.n1501 VSS.n1500 25.6005
R3017 VSS.n1500 VSS.n1497 25.6005
R3018 VSS.n1497 VSS.n1496 25.6005
R3019 VSS.n2012 VSS.n787 25.6005
R3020 VSS.n2012 VSS.n2011 25.6005
R3021 VSS.n2011 VSS.n2010 25.6005
R3022 VSS.n2010 VSS.n2008 25.6005
R3023 VSS.n2008 VSS.n2005 25.6005
R3024 VSS.n2005 VSS.n2004 25.6005
R3025 VSS.n2004 VSS.n2001 25.6005
R3026 VSS.n2001 VSS.n2000 25.6005
R3027 VSS.n2000 VSS.n1997 25.6005
R3028 VSS.n1997 VSS.n1996 25.6005
R3029 VSS.n1996 VSS.n1993 25.6005
R3030 VSS.n1993 VSS.n1992 25.6005
R3031 VSS.n1992 VSS.n1989 25.6005
R3032 VSS.n1989 VSS.n1988 25.6005
R3033 VSS.n1988 VSS.n1985 25.6005
R3034 VSS.n1985 VSS.n1984 25.6005
R3035 VSS.n1984 VSS.n1981 25.6005
R3036 VSS.n1981 VSS.n1980 25.6005
R3037 VSS.n1980 VSS.n1978 25.6005
R3038 VSS.n1978 VSS.n1977 25.6005
R3039 VSS.n1977 VSS.n800 25.6005
R3040 VSS.n1972 VSS.n800 25.6005
R3041 VSS.n1971 VSS.n1970 25.6005
R3042 VSS.n1970 VSS.n1967 25.6005
R3043 VSS.n1967 VSS.n1966 25.6005
R3044 VSS.n1966 VSS.n1963 25.6005
R3045 VSS.n1963 VSS.n1962 25.6005
R3046 VSS.n1962 VSS.n1959 25.6005
R3047 VSS.n1959 VSS.n1958 25.6005
R3048 VSS.n1958 VSS.n1955 25.6005
R3049 VSS.n1955 VSS.n1954 25.6005
R3050 VSS.n1954 VSS.n1951 25.6005
R3051 VSS.n1951 VSS.n1950 25.6005
R3052 VSS.n1950 VSS.n1947 25.6005
R3053 VSS.n1947 VSS.n1946 25.6005
R3054 VSS.n1946 VSS.n1943 25.6005
R3055 VSS.n1943 VSS.n1942 25.6005
R3056 VSS.n1942 VSS.n1939 25.6005
R3057 VSS.n1939 VSS.n1938 25.6005
R3058 VSS.n1938 VSS.n1935 25.6005
R3059 VSS.n1935 VSS.n1934 25.6005
R3060 VSS.n1934 VSS.n1931 25.6005
R3061 VSS.n1931 VSS.n1930 25.6005
R3062 VSS.n1930 VSS.n1927 25.6005
R3063 VSS.n1927 VSS.n1926 25.6005
R3064 VSS.n1923 VSS.n1922 25.6005
R3065 VSS.n1922 VSS.n1919 25.6005
R3066 VSS.n1919 VSS.n1918 25.6005
R3067 VSS.n1918 VSS.n1915 25.6005
R3068 VSS.n1915 VSS.n1914 25.6005
R3069 VSS.n1914 VSS.n1911 25.6005
R3070 VSS.n1911 VSS.n1910 25.6005
R3071 VSS.n1910 VSS.n1907 25.6005
R3072 VSS.n1907 VSS.n1906 25.6005
R3073 VSS.n1906 VSS.n1903 25.6005
R3074 VSS.n1903 VSS.n1902 25.6005
R3075 VSS.n1902 VSS.n1899 25.6005
R3076 VSS.n1899 VSS.n1898 25.6005
R3077 VSS.n1898 VSS.n1895 25.6005
R3078 VSS.n1895 VSS.n1894 25.6005
R3079 VSS.n1894 VSS.n1891 25.6005
R3080 VSS.n1891 VSS.n1890 25.6005
R3081 VSS.n1890 VSS.n1887 25.6005
R3082 VSS.n1887 VSS.n1886 25.6005
R3083 VSS.n1886 VSS.n1883 25.6005
R3084 VSS.n1883 VSS.n1882 25.6005
R3085 VSS.n1882 VSS.n1879 25.6005
R3086 VSS.n1879 VSS.n1878 25.6005
R3087 VSS.n1875 VSS.n1874 25.6005
R3088 VSS.n1874 VSS.n1871 25.6005
R3089 VSS.n1871 VSS.n1870 25.6005
R3090 VSS.n1870 VSS.n1867 25.6005
R3091 VSS.n1867 VSS.n1866 25.6005
R3092 VSS.n1866 VSS.n1863 25.6005
R3093 VSS.n1863 VSS.n1862 25.6005
R3094 VSS.n1862 VSS.n1859 25.6005
R3095 VSS.n1859 VSS.n1858 25.6005
R3096 VSS.n1858 VSS.n1855 25.6005
R3097 VSS.n1855 VSS.n1854 25.6005
R3098 VSS.n1854 VSS.n1851 25.6005
R3099 VSS.n1851 VSS.n1850 25.6005
R3100 VSS.n1850 VSS.n1847 25.6005
R3101 VSS.n1847 VSS.n1846 25.6005
R3102 VSS.n1846 VSS.n1843 25.6005
R3103 VSS.n1843 VSS.n1842 25.6005
R3104 VSS.n1842 VSS.n1839 25.6005
R3105 VSS.n1839 VSS.n1838 25.6005
R3106 VSS.n1838 VSS.n1835 25.6005
R3107 VSS.n1835 VSS.n1834 25.6005
R3108 VSS.n1834 VSS.n1832 25.6005
R3109 VSS.n1390 VSS.n1389 25.6005
R3110 VSS.n1389 VSS.n1388 25.6005
R3111 VSS.n1388 VSS.n1377 25.6005
R3112 VSS.n1380 VSS.n1377 25.6005
R3113 VSS.n1380 VSS.n1379 25.6005
R3114 VSS.n1379 VSS.n1127 25.6005
R3115 VSS.n1487 VSS.n1127 25.6005
R3116 VSS.n1488 VSS.n1487 25.6005
R3117 VSS.n1490 VSS.n1488 25.6005
R3118 VSS.n1490 VSS.n1489 25.6005
R3119 VSS.n1489 VSS.n1104 25.6005
R3120 VSS.n1544 VSS.n1104 25.6005
R3121 VSS.n1545 VSS.n1544 25.6005
R3122 VSS.n1547 VSS.n1545 25.6005
R3123 VSS.n1547 VSS.n1546 25.6005
R3124 VSS.n1568 VSS.n1033 25.6005
R3125 VSS.n1584 VSS.n930 25.6005
R3126 VSS.n1584 VSS.n1583 25.6005
R3127 VSS.n1583 VSS.n1582 25.6005
R3128 VSS.n1615 VSS.n908 25.6005
R3129 VSS.n1616 VSS.n1615 25.6005
R3130 VSS.n1617 VSS.n1616 25.6005
R3131 VSS.n1617 VSS.n886 25.6005
R3132 VSS.n1670 VSS.n886 25.6005
R3133 VSS.n1671 VSS.n1670 25.6005
R3134 VSS.n1672 VSS.n1671 25.6005
R3135 VSS.n1672 VSS.n882 25.6005
R3136 VSS.n1741 VSS.n882 25.6005
R3137 VSS.n1742 VSS.n1741 25.6005
R3138 VSS.n1746 VSS.n1742 25.6005
R3139 VSS.n1746 VSS.n1745 25.6005
R3140 VSS.n1745 VSS.n1744 25.6005
R3141 VSS.n1744 VSS.n843 25.6005
R3142 VSS.n1831 VSS.n843 25.6005
R3143 VSS.n1192 VSS.n649 25.6005
R3144 VSS.n1195 VSS.n1192 25.6005
R3145 VSS.n1196 VSS.n1195 25.6005
R3146 VSS.n1199 VSS.n1196 25.6005
R3147 VSS.n1200 VSS.n1199 25.6005
R3148 VSS.n1203 VSS.n1200 25.6005
R3149 VSS.n1204 VSS.n1203 25.6005
R3150 VSS.n1207 VSS.n1204 25.6005
R3151 VSS.n1208 VSS.n1207 25.6005
R3152 VSS.n1211 VSS.n1208 25.6005
R3153 VSS.n1212 VSS.n1211 25.6005
R3154 VSS.n1215 VSS.n1212 25.6005
R3155 VSS.n1216 VSS.n1215 25.6005
R3156 VSS.n1219 VSS.n1216 25.6005
R3157 VSS.n1220 VSS.n1219 25.6005
R3158 VSS.n1223 VSS.n1220 25.6005
R3159 VSS.n1224 VSS.n1223 25.6005
R3160 VSS.n1227 VSS.n1224 25.6005
R3161 VSS.n1228 VSS.n1227 25.6005
R3162 VSS.n1231 VSS.n1228 25.6005
R3163 VSS.n1232 VSS.n1231 25.6005
R3164 VSS.n1235 VSS.n1232 25.6005
R3165 VSS.n1239 VSS.n1236 25.6005
R3166 VSS.n1240 VSS.n1239 25.6005
R3167 VSS.n1243 VSS.n1240 25.6005
R3168 VSS.n1244 VSS.n1243 25.6005
R3169 VSS.n1247 VSS.n1244 25.6005
R3170 VSS.n1248 VSS.n1247 25.6005
R3171 VSS.n1251 VSS.n1248 25.6005
R3172 VSS.n1252 VSS.n1251 25.6005
R3173 VSS.n1255 VSS.n1252 25.6005
R3174 VSS.n1256 VSS.n1255 25.6005
R3175 VSS.n1259 VSS.n1256 25.6005
R3176 VSS.n1260 VSS.n1259 25.6005
R3177 VSS.n1263 VSS.n1260 25.6005
R3178 VSS.n1264 VSS.n1263 25.6005
R3179 VSS.n1267 VSS.n1264 25.6005
R3180 VSS.n1268 VSS.n1267 25.6005
R3181 VSS.n1271 VSS.n1268 25.6005
R3182 VSS.n1272 VSS.n1271 25.6005
R3183 VSS.n1275 VSS.n1272 25.6005
R3184 VSS.n1276 VSS.n1275 25.6005
R3185 VSS.n1279 VSS.n1276 25.6005
R3186 VSS.n1280 VSS.n1279 25.6005
R3187 VSS.n1283 VSS.n1280 25.6005
R3188 VSS.n1287 VSS.n1284 25.6005
R3189 VSS.n1288 VSS.n1287 25.6005
R3190 VSS.n1291 VSS.n1288 25.6005
R3191 VSS.n1292 VSS.n1291 25.6005
R3192 VSS.n1295 VSS.n1292 25.6005
R3193 VSS.n1296 VSS.n1295 25.6005
R3194 VSS.n1299 VSS.n1296 25.6005
R3195 VSS.n1300 VSS.n1299 25.6005
R3196 VSS.n1303 VSS.n1300 25.6005
R3197 VSS.n1304 VSS.n1303 25.6005
R3198 VSS.n1307 VSS.n1304 25.6005
R3199 VSS.n1308 VSS.n1307 25.6005
R3200 VSS.n1311 VSS.n1308 25.6005
R3201 VSS.n1312 VSS.n1311 25.6005
R3202 VSS.n1315 VSS.n1312 25.6005
R3203 VSS.n1316 VSS.n1315 25.6005
R3204 VSS.n1319 VSS.n1316 25.6005
R3205 VSS.n1320 VSS.n1319 25.6005
R3206 VSS.n1323 VSS.n1320 25.6005
R3207 VSS.n1324 VSS.n1323 25.6005
R3208 VSS.n1327 VSS.n1324 25.6005
R3209 VSS.n1328 VSS.n1327 25.6005
R3210 VSS.n1331 VSS.n1328 25.6005
R3211 VSS.n1335 VSS.n1332 25.6005
R3212 VSS.n1336 VSS.n1335 25.6005
R3213 VSS.n1339 VSS.n1336 25.6005
R3214 VSS.n1340 VSS.n1339 25.6005
R3215 VSS.n1343 VSS.n1340 25.6005
R3216 VSS.n1344 VSS.n1343 25.6005
R3217 VSS.n1347 VSS.n1344 25.6005
R3218 VSS.n1348 VSS.n1347 25.6005
R3219 VSS.n1351 VSS.n1348 25.6005
R3220 VSS.n1352 VSS.n1351 25.6005
R3221 VSS.n1355 VSS.n1352 25.6005
R3222 VSS.n1356 VSS.n1355 25.6005
R3223 VSS.n1359 VSS.n1356 25.6005
R3224 VSS.n1360 VSS.n1359 25.6005
R3225 VSS.n1363 VSS.n1360 25.6005
R3226 VSS.n1364 VSS.n1363 25.6005
R3227 VSS.n1367 VSS.n1364 25.6005
R3228 VSS.n1368 VSS.n1367 25.6005
R3229 VSS.n1369 VSS.n1368 25.6005
R3230 VSS.n1369 VSS.n1154 25.6005
R3231 VSS.n1375 VSS.n1154 25.6005
R3232 VSS.n1376 VSS.n1375 25.6005
R3233 VSS.n2091 VSS.n2090 25.6005
R3234 VSS.n2090 VSS.n2089 25.6005
R3235 VSS.n2089 VSS.n650 25.6005
R3236 VSS.n2083 VSS.n650 25.6005
R3237 VSS.n2083 VSS.n2082 25.6005
R3238 VSS.n2082 VSS.n2081 25.6005
R3239 VSS.n2081 VSS.n654 25.6005
R3240 VSS.n2075 VSS.n654 25.6005
R3241 VSS.n2075 VSS.n2074 25.6005
R3242 VSS.n2074 VSS.n2073 25.6005
R3243 VSS.n2073 VSS.n658 25.6005
R3244 VSS.n2067 VSS.n658 25.6005
R3245 VSS.n2067 VSS.n2066 25.6005
R3246 VSS.n2066 VSS.n2065 25.6005
R3247 VSS.n2065 VSS.n662 25.6005
R3248 VSS.n2059 VSS.n2058 25.6005
R3249 VSS.n1040 VSS.n667 25.6005
R3250 VSS.n1040 VSS.n1039 25.6005
R3251 VSS.n1039 VSS.n769 25.6005
R3252 VSS.n2044 VSS.n774 25.6005
R3253 VSS.n2044 VSS.n2043 25.6005
R3254 VSS.n2043 VSS.n2042 25.6005
R3255 VSS.n2042 VSS.n775 25.6005
R3256 VSS.n2036 VSS.n775 25.6005
R3257 VSS.n2036 VSS.n2035 25.6005
R3258 VSS.n2035 VSS.n2034 25.6005
R3259 VSS.n2034 VSS.n779 25.6005
R3260 VSS.n2028 VSS.n779 25.6005
R3261 VSS.n2028 VSS.n2027 25.6005
R3262 VSS.n2027 VSS.n2026 25.6005
R3263 VSS.n2026 VSS.n783 25.6005
R3264 VSS.n2020 VSS.n783 25.6005
R3265 VSS.n2020 VSS.n2019 25.6005
R3266 VSS.n2019 VSS.n2018 25.6005
R3267 VSS.n1751 VSS.n875 25.6005
R3268 VSS.n1752 VSS.n1751 25.6005
R3269 VSS.n1753 VSS.n1752 25.6005
R3270 VSS.n1753 VSS.n849 25.6005
R3271 VSS.n1826 VSS.n849 25.6005
R3272 VSS.n1826 VSS.n1825 25.6005
R3273 VSS.n1825 VSS.n1824 25.6005
R3274 VSS.n1824 VSS.n1823 25.6005
R3275 VSS.n1823 VSS.n850 25.6005
R3276 VSS.n857 VSS.n850 25.6005
R3277 VSS.n1816 VSS.n857 25.6005
R3278 VSS.n1735 VSS.n1734 25.6005
R3279 VSS.n1734 VSS.n1733 25.6005
R3280 VSS.n1733 VSS.n1730 25.6005
R3281 VSS.n1730 VSS.n1729 25.6005
R3282 VSS.n1729 VSS.n1726 25.6005
R3283 VSS.n1726 VSS.n1725 25.6005
R3284 VSS.n1725 VSS.n1722 25.6005
R3285 VSS.n1722 VSS.n1721 25.6005
R3286 VSS.n1721 VSS.n1718 25.6005
R3287 VSS.n1718 VSS.n1717 25.6005
R3288 VSS.n1717 VSS.n1714 25.6005
R3289 VSS.n1714 VSS.n1713 25.6005
R3290 VSS.n1713 VSS.n1710 25.6005
R3291 VSS.n1710 VSS.n1709 25.6005
R3292 VSS.n1709 VSS.n1706 25.6005
R3293 VSS.n1706 VSS.n1705 25.6005
R3294 VSS.n1705 VSS.n1702 25.6005
R3295 VSS.n1702 VSS.n1701 25.6005
R3296 VSS.n1701 VSS.n1698 25.6005
R3297 VSS.n1698 VSS.n1697 25.6005
R3298 VSS.n1697 VSS.n1694 25.6005
R3299 VSS.n1694 VSS.n1693 25.6005
R3300 VSS.n1689 VSS.n1688 25.6005
R3301 VSS.n1688 VSS.n1687 25.6005
R3302 VSS.n1687 VSS.n870 25.6005
R3303 VSS.n1759 VSS.n870 25.6005
R3304 VSS.n1760 VSS.n1759 25.6005
R3305 VSS.n1762 VSS.n1760 25.6005
R3306 VSS.n1763 VSS.n1762 25.6005
R3307 VSS.n1765 VSS.n1763 25.6005
R3308 VSS.n1766 VSS.n1765 25.6005
R3309 VSS.n1767 VSS.n1766 25.6005
R3310 VSS.n1768 VSS.n1767 25.6005
R3311 VSS.n1815 VSS.n1814 25.6005
R3312 VSS.n1814 VSS.n858 25.6005
R3313 VSS.n1809 VSS.n858 25.6005
R3314 VSS.n1809 VSS.n1808 25.6005
R3315 VSS.n1808 VSS.n860 25.6005
R3316 VSS.n1803 VSS.n860 25.6005
R3317 VSS.n1803 VSS.n1802 25.6005
R3318 VSS.n1802 VSS.n1801 25.6005
R3319 VSS.n1801 VSS.n862 25.6005
R3320 VSS.n1792 VSS.n1791 25.6005
R3321 VSS.n1791 VSS.n865 25.6005
R3322 VSS.n1785 VSS.n865 25.6005
R3323 VSS.n1785 VSS.n1784 25.6005
R3324 VSS.n1784 VSS.n1783 25.6005
R3325 VSS.n1783 VSS.n867 25.6005
R3326 VSS.n1777 VSS.n867 25.6005
R3327 VSS.n1777 VSS.n1776 25.6005
R3328 VSS.n1776 VSS.n1775 25.6005
R3329 VSS.n1775 VSS.n869 25.6005
R3330 VSS.n1769 VSS.n869 25.6005
R3331 VSS.n542 VSS.n537 25.6005
R3332 VSS.n542 VSS.n541 25.6005
R3333 VSS.n548 VSS.n541 25.6005
R3334 VSS.n549 VSS.n548 25.6005
R3335 VSS.n555 VSS.n554 25.6005
R3336 VSS.n556 VSS.n555 25.6005
R3337 VSS.n556 VSS.n529 25.6005
R3338 VSS.n567 VSS.n529 25.6005
R3339 VSS.n568 VSS.n567 25.6005
R3340 VSS.n569 VSS.n568 25.6005
R3341 VSS.n569 VSS.n440 25.6005
R3342 VSS.n2193 VSS.n440 25.6005
R3343 VSS.n2193 VSS.n2192 25.6005
R3344 VSS.n2192 VSS.n2191 25.6005
R3345 VSS.n2191 VSS.n441 25.6005
R3346 VSS.n2185 VSS.n441 25.6005
R3347 VSS.n2185 VSS.n2184 25.6005
R3348 VSS.n2184 VSS.n2183 25.6005
R3349 VSS.n2183 VSS.n448 25.6005
R3350 VSS.n2177 VSS.n448 25.6005
R3351 VSS.n2177 VSS.n2176 25.6005
R3352 VSS.n2176 VSS.n2175 25.6005
R3353 VSS.n2175 VSS.n455 25.6005
R3354 VSS.n2169 VSS.n455 25.6005
R3355 VSS.n2169 VSS.n2168 25.6005
R3356 VSS.n2168 VSS.n2167 25.6005
R3357 VSS.n2167 VSS.n462 25.6005
R3358 VSS.n2161 VSS.n462 25.6005
R3359 VSS.n2161 VSS.n2160 25.6005
R3360 VSS.n2160 VSS.n2159 25.6005
R3361 VSS.n2159 VSS.n469 25.6005
R3362 VSS.n2153 VSS.n469 25.6005
R3363 VSS.n2153 VSS.n2152 25.6005
R3364 VSS.n2152 VSS.n2151 25.6005
R3365 VSS.n2151 VSS.n476 25.6005
R3366 VSS.n2145 VSS.n476 25.6005
R3367 VSS.n2145 VSS.n2144 25.6005
R3368 VSS.n2144 VSS.n2143 25.6005
R3369 VSS.n2143 VSS.n483 25.6005
R3370 VSS.n2137 VSS.n483 25.6005
R3371 VSS.n2137 VSS.n2136 25.6005
R3372 VSS.n2136 VSS.n2135 25.6005
R3373 VSS.n2135 VSS.n490 25.6005
R3374 VSS.n2129 VSS.n490 25.6005
R3375 VSS.n2129 VSS.n2128 25.6005
R3376 VSS.n2128 VSS.n2127 25.6005
R3377 VSS.n2127 VSS.n497 25.6005
R3378 VSS.n2121 VSS.n497 25.6005
R3379 VSS.n2121 VSS.n2120 25.6005
R3380 VSS.n2120 VSS.n2119 25.6005
R3381 VSS.n2119 VSS.n504 25.6005
R3382 VSS.n2113 VSS.n504 25.6005
R3383 VSS.n2113 VSS.n2112 25.6005
R3384 VSS.n2112 VSS.n2111 25.6005
R3385 VSS.n2111 VSS.n511 25.6005
R3386 VSS.n2105 VSS.n511 25.6005
R3387 VSS.n2105 VSS.n2104 25.6005
R3388 VSS.n2099 VSS.n520 25.6005
R3389 VSS.n524 VSS.n520 25.6005
R3390 VSS.n633 VSS.n524 25.6005
R3391 VSS.n550 VSS.n533 25.6005
R3392 VSS.n560 VSS.n533 25.6005
R3393 VSS.n561 VSS.n560 25.6005
R3394 VSS.n563 VSS.n561 25.6005
R3395 VSS.n563 VSS.n562 25.6005
R3396 VSS.n562 VSS.n525 25.6005
R3397 VSS.n574 VSS.n525 25.6005
R3398 VSS.n575 VSS.n574 25.6005
R3399 VSS.n577 VSS.n575 25.6005
R3400 VSS.n578 VSS.n577 25.6005
R3401 VSS.n579 VSS.n578 25.6005
R3402 VSS.n580 VSS.n579 25.6005
R3403 VSS.n582 VSS.n580 25.6005
R3404 VSS.n583 VSS.n582 25.6005
R3405 VSS.n584 VSS.n583 25.6005
R3406 VSS.n585 VSS.n584 25.6005
R3407 VSS.n587 VSS.n585 25.6005
R3408 VSS.n588 VSS.n587 25.6005
R3409 VSS.n589 VSS.n588 25.6005
R3410 VSS.n590 VSS.n589 25.6005
R3411 VSS.n592 VSS.n590 25.6005
R3412 VSS.n593 VSS.n592 25.6005
R3413 VSS.n594 VSS.n593 25.6005
R3414 VSS.n595 VSS.n594 25.6005
R3415 VSS.n597 VSS.n595 25.6005
R3416 VSS.n598 VSS.n597 25.6005
R3417 VSS.n600 VSS.n598 25.6005
R3418 VSS.n601 VSS.n600 25.6005
R3419 VSS.n603 VSS.n601 25.6005
R3420 VSS.n604 VSS.n603 25.6005
R3421 VSS.n605 VSS.n604 25.6005
R3422 VSS.n606 VSS.n605 25.6005
R3423 VSS.n608 VSS.n606 25.6005
R3424 VSS.n609 VSS.n608 25.6005
R3425 VSS.n610 VSS.n609 25.6005
R3426 VSS.n611 VSS.n610 25.6005
R3427 VSS.n613 VSS.n611 25.6005
R3428 VSS.n614 VSS.n613 25.6005
R3429 VSS.n615 VSS.n614 25.6005
R3430 VSS.n616 VSS.n615 25.6005
R3431 VSS.n618 VSS.n616 25.6005
R3432 VSS.n619 VSS.n618 25.6005
R3433 VSS.n620 VSS.n619 25.6005
R3434 VSS.n621 VSS.n620 25.6005
R3435 VSS.n623 VSS.n621 25.6005
R3436 VSS.n624 VSS.n623 25.6005
R3437 VSS.n625 VSS.n624 25.6005
R3438 VSS.n626 VSS.n625 25.6005
R3439 VSS.n628 VSS.n626 25.6005
R3440 VSS.n629 VSS.n628 25.6005
R3441 VSS.n630 VSS.n629 25.6005
R3442 VSS.n631 VSS.n630 25.6005
R3443 VSS.n632 VSS.n631 25.6005
R3444 VSS.n1554 VSS.n1553 25.6005
R3445 VSS.n1553 VSS.n1052 25.6005
R3446 VSS.n1064 VSS.n1052 25.6005
R3447 VSS.n1067 VSS.n1064 25.6005
R3448 VSS.n1068 VSS.n1067 25.6005
R3449 VSS.n1071 VSS.n1068 25.6005
R3450 VSS.n1072 VSS.n1071 25.6005
R3451 VSS.n1075 VSS.n1072 25.6005
R3452 VSS.n1076 VSS.n1075 25.6005
R3453 VSS.n1079 VSS.n1076 25.6005
R3454 VSS.n1080 VSS.n1079 25.6005
R3455 VSS.n1083 VSS.n1080 25.6005
R3456 VSS.n1084 VSS.n1083 25.6005
R3457 VSS.n1087 VSS.n1084 25.6005
R3458 VSS.n1088 VSS.n1087 25.6005
R3459 VSS.n1091 VSS.n1088 25.6005
R3460 VSS.n1092 VSS.n1091 25.6005
R3461 VSS.n1095 VSS.n1092 25.6005
R3462 VSS.n1097 VSS.n1095 25.6005
R3463 VSS.n1098 VSS.n1097 25.6005
R3464 VSS.n1099 VSS.n1098 25.6005
R3465 VSS.n1099 VSS.n1045 25.6005
R3466 VSS.n1556 VSS.n1555 25.6005
R3467 VSS.n1555 VSS.n923 25.6005
R3468 VSS.n1589 VSS.n923 25.6005
R3469 VSS.n1590 VSS.n1589 25.6005
R3470 VSS.n1591 VSS.n1590 25.6005
R3471 VSS.n1591 VSS.n914 25.6005
R3472 VSS.n1607 VSS.n914 25.6005
R3473 VSS.n1608 VSS.n1607 25.6005
R3474 VSS.n1610 VSS.n1608 25.6005
R3475 VSS.n1610 VSS.n1609 25.6005
R3476 VSS.n1609 VSS.n902 25.6005
R3477 VSS.n1664 VSS.n1663 25.6005
R3478 VSS.n1663 VSS.n1662 25.6005
R3479 VSS.n1662 VSS.n1661 25.6005
R3480 VSS.n1661 VSS.n1659 25.6005
R3481 VSS.n1659 VSS.n1656 25.6005
R3482 VSS.n1656 VSS.n1655 25.6005
R3483 VSS.n1655 VSS.n1652 25.6005
R3484 VSS.n1652 VSS.n1651 25.6005
R3485 VSS.n1651 VSS.n1648 25.6005
R3486 VSS.n1648 VSS.n1647 25.6005
R3487 VSS.n1647 VSS.n1644 25.6005
R3488 VSS.n1644 VSS.n1643 25.6005
R3489 VSS.n1643 VSS.n1640 25.6005
R3490 VSS.n1640 VSS.n1639 25.6005
R3491 VSS.n1639 VSS.n1636 25.6005
R3492 VSS.n1636 VSS.n1635 25.6005
R3493 VSS.n1635 VSS.n1632 25.6005
R3494 VSS.n1632 VSS.n1631 25.6005
R3495 VSS.n1631 VSS.n1628 25.6005
R3496 VSS.n1628 VSS.n1627 25.6005
R3497 VSS.n1627 VSS.n1624 25.6005
R3498 VSS.n1624 VSS.n1623 25.6005
R3499 VSS.n1561 VSS.n1560 25.6005
R3500 VSS.n1563 VSS.n1561 25.6005
R3501 VSS.n1563 VSS.n1562 25.6005
R3502 VSS.n1562 VSS.n919 25.6005
R3503 VSS.n1595 VSS.n919 25.6005
R3504 VSS.n1596 VSS.n1595 25.6005
R3505 VSS.n1602 VSS.n1596 25.6005
R3506 VSS.n1598 VSS.n1597 25.6005
R3507 VSS.n1597 VSS.n903 25.6005
R3508 VSS.t112 VSS.n1819 25.0064
R3509 VSS.n2197 VSS.n2195 24.8841
R3510 VSS.n302 VSS.n296 24.8476
R3511 VSS.n357 VSS.n351 24.8476
R3512 VSS.n65 VSS.n47 24.8476
R3513 VSS.n19 VSS.n18 24.8476
R3514 VSS.n285 VSS.n230 24.8476
R3515 VSS.n2408 VSS.n2407 24.8476
R3516 VSS.n1470 VSS.n1121 24.8476
R3517 VSS.n752 VSS.n751 24.8476
R3518 VSS.n691 VSS.n687 24.8476
R3519 VSS.n1014 VSS.n984 24.8476
R3520 VSS.n953 VSS.n950 24.8476
R3521 VSS.n1577 VSS.n1031 24.8476
R3522 VSS.n2051 VSS.n2050 24.8476
R3523 VSS.n60 VSS.n59 24.75
R3524 VSS.n23 VSS.n22 24.75
R3525 VSS.n315 VSS.n291 24.2609
R3526 VSS.n309 VSS.n289 24.2609
R3527 VSS.n370 VSS.n364 24.2609
R3528 VSS.n375 VSS.n366 24.2609
R3529 VSS.n53 VSS.n49 24.2609
R3530 VSS.n27 VSS.n6 24.2609
R3531 VSS.n2103 VSS.n518 23.7181
R3532 VSS.n1542 VSS.n1540 23.4436
R3533 VSS.n315 VSS.n292 23.3417
R3534 VSS.n309 VSS.n290 23.3417
R3535 VSS.n299 VSS.n295 23.3417
R3536 VSS.n370 VSS.n365 23.3417
R3537 VSS.n375 VSS.n367 23.3417
R3538 VSS.n354 VSS.n350 23.3417
R3539 VSS.n69 VSS.n68 23.3417
R3540 VSS.n53 VSS.n50 23.3417
R3541 VSS.n28 VSS.n27 23.3417
R3542 VSS.n15 VSS.n10 23.3417
R3543 VSS.n748 VSS.n722 23.3417
R3544 VSS.n692 VSS.n685 23.3417
R3545 VSS.n1013 VSS.n986 23.3417
R3546 VSS.n957 VSS.n956 23.3417
R3547 VSS.n1749 VSS.n877 22.9226
R3548 VSS.n1755 VSS.n872 22.9226
R3549 VSS.n1828 VSS.n845 22.9226
R3550 VSS.n1546 VSS.n1032 22.5887
R3551 VSS.n666 VSS.n662 22.5887
R3552 VSS.n303 VSS.n302 22.4252
R3553 VSS.n358 VSS.n357 22.4252
R3554 VSS.n2210 VSS.t120 22.4016
R3555 VSS.n2346 VSS.t17 22.4016
R3556 VSS.n1569 VSS.n930 22.2123
R3557 VSS.n2057 VSS.n667 22.2123
R3558 VSS.n319 VSS.n318 21.8358
R3559 VSS.n322 VSS.n288 21.8358
R3560 VSS.n305 VSS.n294 21.8358
R3561 VSS.n382 VSS.n363 21.8358
R3562 VSS.n379 VSS.n378 21.8358
R3563 VSS.n360 VSS.n349 21.8358
R3564 VSS.n71 VSS.n45 21.8358
R3565 VSS.n57 VSS.n56 21.8358
R3566 VSS.n30 VSS.n5 21.8358
R3567 VSS.n14 VSS.n11 21.8358
R3568 VSS.n1474 VSS.n1473 21.8358
R3569 VSS.n747 VSS.n724 21.8358
R3570 VSS.n696 VSS.n695 21.8358
R3571 VSS.n1010 VSS.n1009 21.8358
R3572 VSS.n960 VSS.n948 21.8358
R3573 VSS.n2274 VSS.t0 21.3597
R3574 VSS.t113 VSS.n157 21.3597
R3575 VSS.n388 VSS.n230 21.0829
R3576 VSS.n2407 VSS.n2405 21.0829
R3577 VSS.n1035 VSS.n664 20.4928
R3578 VSS.n744 VSS.n743 20.3299
R3579 VSS.n699 VSS.n683 20.3299
R3580 VSS.n1006 VSS.n988 20.3299
R3581 VSS.n961 VSS.n946 20.3299
R3582 VSS.n2230 VSS.t23 20.3178
R3583 VSS.n133 VSS.t107 20.3178
R3584 VSS.n1757 VSS.t19 20.3178
R3585 VSS.n278 VSS.n231 19.9534
R3586 VSS.n2411 VSS.n2410 19.9534
R3587 VSS.n1558 VSS.n1047 19.7969
R3588 VSS.n1050 VSS.n1048 19.7969
R3589 VSS.n1587 VSS.n925 19.7969
R3590 VSS.n1586 VSS.n927 19.7969
R3591 VSS.n1593 VSS.n921 19.7969
R3592 VSS.n1605 VSS.n916 19.7969
R3593 VSS.n1604 VSS.n910 19.7969
R3594 VSS.n1613 VSS.n1612 19.7969
R3595 VSS.n906 VSS.n905 19.7969
R3596 VSS.n1620 VSS.n1619 19.7969
R3597 VSS.n740 VSS.n726 18.824
R3598 VSS.n700 VSS.n681 18.824
R3599 VSS.n1005 VSS.n990 18.824
R3600 VSS.n965 VSS.n964 18.824
R3601 VSS.n1454 VSS.n1392 18.7549
R3602 VSS.n1151 VSS.n1146 18.7549
R3603 VSS.n1385 VSS.n1142 18.7549
R3604 VSS.n1381 VSS.n1137 18.7549
R3605 VSS.n1485 VSS.n1130 18.7549
R3606 VSS.n1492 VSS.n1123 18.7549
R3607 VSS.n1576 VSS.n908 18.4476
R3608 VSS.n774 VSS.n768 18.4476
R3609 VSS.n884 VSS.t2 18.234
R3610 VSS.n1795 VSS.n864 18.0711
R3611 VSS.n1600 VSS.n1599 18.0711
R3612 VSS.n1466 VSS.t30 17.713
R3613 VSS.t110 VSS.n1579 17.713
R3614 VSS.t14 VSS.n802 17.713
R3615 VSS.n739 VSS.n728 17.3181
R3616 VSS.n705 VSS.n704 17.3181
R3617 VSS.n1002 VSS.n1001 17.3181
R3618 VSS.n968 VSS.n944 17.3181
R3619 VSS.n732 VSS.n731 17.1928
R3620 VSS.n711 VSS.n710 17.1928
R3621 VSS.n995 VSS.n994 17.1928
R3622 VSS.n973 VSS.n940 17.1928
R3623 VSS.n1125 VSS.t10 17.1921
R3624 VSS.n1460 VSS.n1146 16.6711
R3625 VSS.n1386 VSS.n1385 16.6711
R3626 VSS.n1466 VSS.n1142 16.6711
R3627 VSS.n1382 VSS.n1381 16.6711
R3628 VSS.n1477 VSS.n1137 16.6711
R3629 VSS.n1130 VSS.n1129 16.6711
R3630 VSS.n1485 VSS.n1484 16.6711
R3631 VSS.n1132 VSS.n1123 16.6711
R3632 VSS.n1493 VSS.n1492 16.6711
R3633 VSS.n1460 VSS.t36 16.1502
R3634 VSS.n736 VSS.n735 15.8123
R3635 VSS.n708 VSS.n679 15.8123
R3636 VSS.n998 VSS.n992 15.8123
R3637 VSS.n969 VSS.n942 15.8123
R3638 VSS.n1558 VSS.n1048 15.6292
R3639 VSS.n1565 VSS.n925 15.6292
R3640 VSS.n1587 VSS.n1586 15.6292
R3641 VSS.n927 VSS.n921 15.6292
R3642 VSS.n1579 VSS.n916 15.6292
R3643 VSS.n1605 VSS.n1604 15.6292
R3644 VSS.n1613 VSS.n910 15.6292
R3645 VSS.n1619 VSS.n905 15.6292
R3646 VSS.n1620 VSS.n888 15.6292
R3647 VSS.n2223 VSS.t23 15.1082
R3648 VSS.n2334 VSS.t107 15.1082
R3649 VSS.n1668 VSS.n1667 15.1082
R3650 VSS.n319 VSS.n308 14.5711
R3651 VSS.n323 VSS.n322 14.5711
R3652 VSS.n306 VSS.n305 14.5711
R3653 VSS.n383 VSS.n382 14.5711
R3654 VSS.n379 VSS.n368 14.5711
R3655 VSS.n361 VSS.n360 14.5711
R3656 VSS.n72 VSS.n71 14.5711
R3657 VSS.n57 VSS.n51 14.5711
R3658 VSS.n31 VSS.n30 14.5711
R3659 VSS.n11 VSS.n3 14.5711
R3660 VSS.n732 VSS.n730 14.3064
R3661 VSS.n710 VSS.n709 14.3064
R3662 VSS.n997 VSS.n994 14.3064
R3663 VSS.n973 VSS.n972 14.3064
R3664 VSS.t0 VSS.n165 14.0663
R3665 VSS.n2286 VSS.t113 14.0663
R3666 VSS.n1794 VSS.n1792 13.5534
R3667 VSS.n1602 VSS.n1601 13.5534
R3668 VSS.n1550 VSS.t9 13.5454
R3669 VSS.n2100 VSS.n518 13.177
R3670 VSS.n2217 VSS.t120 13.0244
R3671 VSS.n125 VSS.t17 13.0244
R3672 VSS.n1690 VSS.t12 13.0244
R3673 VSS.n1690 VSS.n877 12.5035
R3674 VSS.n1749 VSS.n1748 12.5035
R3675 VSS.n1748 VSS.t129 12.5035
R3676 VSS.n879 VSS.n872 12.5035
R3677 VSS.n1755 VSS.n873 12.5035
R3678 VSS.n1757 VSS.n845 12.5035
R3679 VSS.n1829 VSS.n1828 12.5035
R3680 VSS.n2100 VSS.n2099 12.424
R3681 VSS.n1795 VSS.n1794 12.0476
R3682 VSS.n1601 VSS.n1600 12.0476
R3683 VSS.n1540 VSS.n1106 11.9825
R3684 VSS.n1593 VSS.t13 11.9825
R3685 VSS.n735 VSS.n730 11.2946
R3686 VSS.n709 VSS.n708 11.2946
R3687 VSS.n998 VSS.n997 11.2946
R3688 VSS.n972 VSS.n942 11.2946
R3689 VSS.n1023 VSS.n1022 11.0636
R3690 VSS.n1024 VSS.n982 11.0636
R3691 VSS.n1025 VSS.n981 11.0636
R3692 VSS.n1026 VSS.n934 11.0636
R3693 VSS.n975 VSS.n939 11.0636
R3694 VSS.n977 VSS.n976 11.0636
R3695 VSS.n979 VSS.n978 11.0636
R3696 VSS.n980 VSS.n933 11.0636
R3697 VSS.n1028 VSS.n1027 11.0636
R3698 VSS.n760 VSS.n759 11.0636
R3699 VSS.n761 VSS.n719 11.0636
R3700 VSS.n762 VSS.n718 11.0636
R3701 VSS.n763 VSS.n671 11.0636
R3702 VSS.n712 VSS.n676 11.0636
R3703 VSS.n714 VSS.n713 11.0636
R3704 VSS.n716 VSS.n715 11.0636
R3705 VSS.n717 VSS.n670 11.0636
R3706 VSS.n765 VSS.n764 11.0636
R3707 VSS.n1541 VSS.t9 10.9406
R3708 VSS.n1550 VSS.n1549 10.9406
R3709 VSS.t127 VSS.n1151 10.4196
R3710 VSS.n1484 VSS.t116 10.4196
R3711 VSS.t126 VSS.n1565 10.4196
R3712 VSS.t129 VSS.n879 10.4196
R3713 VSS.n1820 VSS.t112 10.4196
R3714 VSS.t79 VSS.n1035 10.2467
R3715 VSS.t13 VSS.n772 10.2467
R3716 VSS.n1129 VSS.t39 9.89868
R3717 VSS.n1739 VSS.t12 9.89868
R3718 VSS.n736 VSS.n728 9.78874
R3719 VSS.n705 VSS.n679 9.78874
R3720 VSS.n1001 VSS.n992 9.78874
R3721 VSS.n969 VSS.n968 9.78874
R3722 VSS.n752 VSS.n720 9.58499
R3723 VSS.n689 VSS.n687 9.58499
R3724 VSS.n1016 VSS.n984 9.58499
R3725 VSS.n953 VSS.n952 9.58499
R3726 VSS.n2101 VSS.n520 9.52595
R3727 VSS.n2410 VSS.n2409 9.49023
R3728 VSS.n286 VSS.n231 9.49023
R3729 VSS.n2052 VSS.n768 9.49023
R3730 VSS.n1576 VSS.n1575 9.49023
R3731 VSS.n1570 VSS.n1032 9.49023
R3732 VSS.n2056 VSS.n666 9.49023
R3733 VSS.n1601 VSS.n1 9.36151
R3734 VSS.n1473 VSS.n2 9.36002
R3735 VSS.n1470 VSS.n2 9.36002
R3736 VSS.n1599 VSS.n1 9.35854
R3737 VSS.n310 VSS.n309 9.3005
R3738 VSS.n288 VSS.n287 9.3005
R3739 VSS.n302 VSS.n301 9.3005
R3740 VSS.n300 VSS.n299 9.3005
R3741 VSS.n294 VSS.n293 9.3005
R3742 VSS.n316 VSS.n315 9.3005
R3743 VSS.n318 VSS.n317 9.3005
R3744 VSS.n376 VSS.n375 9.3005
R3745 VSS.n378 VSS.n377 9.3005
R3746 VSS.n357 VSS.n356 9.3005
R3747 VSS.n355 VSS.n354 9.3005
R3748 VSS.n349 VSS.n348 9.3005
R3749 VSS.n371 VSS.n370 9.3005
R3750 VSS.n363 VSS.n362 9.3005
R3751 VSS.n54 VSS.n53 9.3005
R3752 VSS.n56 VSS.n55 9.3005
R3753 VSS.n66 VSS.n65 9.3005
R3754 VSS.n68 VSS.n67 9.3005
R3755 VSS.n45 VSS.n44 9.3005
R3756 VSS.n19 VSS.n9 9.3005
R3757 VSS.n12 VSS.n10 9.3005
R3758 VSS.n14 VSS.n13 9.3005
R3759 VSS.n27 VSS.n26 9.3005
R3760 VSS.n5 VSS.n4 9.3005
R3761 VSS.n388 VSS.n387 9.3005
R3762 VSS.n386 VSS.n228 9.3005
R3763 VSS.n286 VSS.n285 9.3005
R3764 VSS.n2405 VSS.n75 9.3005
R3765 VSS.n2409 VSS.n2408 9.3005
R3766 VSS.n2454 VSS.n2453 9.3005
R3767 VSS.n753 VSS.n752 9.3005
R3768 VSS.n722 VSS.n721 9.3005
R3769 VSS.n747 VSS.n746 9.3005
R3770 VSS.n745 VSS.n744 9.3005
R3771 VSS.n726 VSS.n725 9.3005
R3772 VSS.n739 VSS.n738 9.3005
R3773 VSS.n737 VSS.n736 9.3005
R3774 VSS.n730 VSS.n729 9.3005
R3775 VSS.n687 VSS.n686 9.3005
R3776 VSS.n693 VSS.n692 9.3005
R3777 VSS.n695 VSS.n694 9.3005
R3778 VSS.n683 VSS.n682 9.3005
R3779 VSS.n701 VSS.n700 9.3005
R3780 VSS.n704 VSS.n703 9.3005
R3781 VSS.n702 VSS.n679 9.3005
R3782 VSS.n709 VSS.n678 9.3005
R3783 VSS.n984 VSS.n983 9.3005
R3784 VSS.n1013 VSS.n1012 9.3005
R3785 VSS.n1011 VSS.n1010 9.3005
R3786 VSS.n988 VSS.n987 9.3005
R3787 VSS.n1005 VSS.n1004 9.3005
R3788 VSS.n1003 VSS.n1002 9.3005
R3789 VSS.n992 VSS.n991 9.3005
R3790 VSS.n997 VSS.n996 9.3005
R3791 VSS.n954 VSS.n953 9.3005
R3792 VSS.n956 VSS.n955 9.3005
R3793 VSS.n948 VSS.n947 9.3005
R3794 VSS.n962 VSS.n961 9.3005
R3795 VSS.n964 VSS.n963 9.3005
R3796 VSS.n944 VSS.n943 9.3005
R3797 VSS.n970 VSS.n969 9.3005
R3798 VSS.n972 VSS.n971 9.3005
R3799 VSS.n1575 VSS.n1031 9.3005
R3800 VSS.n1584 VSS.n1030 9.3005
R3801 VSS.n1570 VSS.n1569 9.3005
R3802 VSS.n2052 VSS.n2051 9.3005
R3803 VSS.n2057 VSS.n2056 9.3005
R3804 VSS.n1040 VSS.n767 9.3005
R3805 VSS.n1793 VSS.n864 9.3005
R3806 VSS.n1794 VSS.n1793 9.3005
R3807 VSS.n2101 VSS.n2100 9.3005
R3808 VSS.n2103 VSS.n2102 9.3005
R3809 VSS.n1477 VSS.t39 8.85676
R3810 VSS.t116 VSS.n1132 8.33581
R3811 VSS.n1050 VSS.n664 8.33581
R3812 VSS.n740 VSS.n739 8.28285
R3813 VSS.n704 VSS.n681 8.28285
R3814 VSS.n1002 VSS.n990 8.28285
R3815 VSS.n965 VSS.n944 8.28285
R3816 VSS.n303 VSS.n298 8.2073
R3817 VSS.n358 VSS.n353 8.2073
R3818 VSS.n2236 VSS.t25 7.81485
R3819 VSS.n2322 VSS.t3 7.81485
R3820 VSS.n1738 VSS.n1737 7.81485
R3821 VSS.n864 VSS.n862 7.52991
R3822 VSS.n1599 VSS.n1598 7.52991
R3823 VSS.n2087 VSS.t36 7.3192
R3824 VSS.n2022 VSS.t19 7.3192
R3825 VSS.n1566 VSS.n664 7.29389
R3826 VSS.n1573 VSS.n1572 7.25768
R3827 VSS.n2054 VSS.n519 7.25768
R3828 VSS.n2156 VSS.n472 7.24494
R3829 VSS.n1577 VSS.n1576 7.15344
R3830 VSS.n2050 VSS.n768 7.15344
R3831 VSS.n743 VSS.n726 6.77697
R3832 VSS.n700 VSS.n699 6.77697
R3833 VSS.n1006 VSS.n1005 6.77697
R3834 VSS.n964 VSS.n946 6.77697
R3835 VSS.t5 VSS.n173 6.77294
R3836 VSS.n2298 VSS.t31 6.77294
R3837 VSS.n314 VSS.n291 6.41949
R3838 VSS.n311 VSS.n289 6.41949
R3839 VSS.n372 VSS.n364 6.41949
R3840 VSS.n374 VSS.n366 6.41949
R3841 VSS.n52 VSS.n49 6.41949
R3842 VSS.n25 VSS.n6 6.41949
R3843 VSS.n1392 VSS.t127 6.25198
R3844 VSS.t100 VSS.n320 5.8005
R3845 VSS.n320 VSS.t56 5.8005
R3846 VSS.n321 VSS.t111 5.8005
R3847 VSS.n321 VSS.t100 5.8005
R3848 VSS.n304 VSS.t109 5.8005
R3849 VSS.n304 VSS.t48 5.8005
R3850 VSS.n381 VSS.t67 5.8005
R3851 VSS.n381 VSS.t65 5.8005
R3852 VSS.t65 VSS.n380 5.8005
R3853 VSS.n380 VSS.t123 5.8005
R3854 VSS.n359 VSS.t60 5.8005
R3855 VSS.n359 VSS.t21 5.8005
R3856 VSS.n325 VSS.t135 5.8005
R3857 VSS.n325 VSS.t122 5.8005
R3858 VSS.n329 VSS.t16 5.8005
R3859 VSS.n329 VSS.t7 5.8005
R3860 VSS.n333 VSS.t136 5.8005
R3861 VSS.n333 VSS.t134 5.8005
R3862 VSS.n337 VSS.t8 5.8005
R3863 VSS.n337 VSS.t132 5.8005
R3864 VSS.n341 VSS.t26 5.8005
R3865 VSS.n341 VSS.t131 5.8005
R3866 VSS.n345 VSS.t121 5.8005
R3867 VSS.n345 VSS.t24 5.8005
R3868 VSS.n327 VSS.t4 5.8005
R3869 VSS.n327 VSS.t124 5.8005
R3870 VSS.n331 VSS.t119 5.8005
R3871 VSS.n331 VSS.t118 5.8005
R3872 VSS.n335 VSS.t27 5.8005
R3873 VSS.n335 VSS.t130 5.8005
R3874 VSS.n339 VSS.t138 5.8005
R3875 VSS.n339 VSS.t22 5.8005
R3876 VSS.n343 VSS.t117 5.8005
R3877 VSS.n343 VSS.t115 5.8005
R3878 VSS.n58 VSS.t18 5.8005
R3879 VSS.t63 VSS.n58 5.8005
R3880 VSS.n59 VSS.t63 5.8005
R3881 VSS.n59 VSS.t87 5.8005
R3882 VSS.n41 VSS.t105 5.8005
R3883 VSS.n41 VSS.t108 5.8005
R3884 VSS.n39 VSS.t32 5.8005
R3885 VSS.n39 VSS.t133 5.8005
R3886 VSS.n37 VSS.t1 5.8005
R3887 VSS.n37 VSS.t114 5.8005
R3888 VSS.n35 VSS.t29 5.8005
R3889 VSS.n35 VSS.t6 5.8005
R3890 VSS.n33 VSS.t137 5.8005
R3891 VSS.n33 VSS.t106 5.8005
R3892 VSS.n29 VSS.t96 5.8005
R3893 VSS.n29 VSS.t125 5.8005
R3894 VSS.n22 VSS.t98 5.8005
R3895 VSS.n22 VSS.t96 5.8005
R3896 VSS.n2204 VSS.t20 5.73102
R3897 VSS.n117 VSS.t62 5.73102
R3898 VSS.t79 VSS.t126 5.73102
R3899 VSS.t11 VSS.t51 5.73102
R3900 VSS.n232 VSS.n231 5.64756
R3901 VSS.n2410 VSS.n2401 5.64756
R3902 VSS.n66 VSS.n62 5.37662
R3903 VSS.n21 VSS.n9 5.37662
R3904 VSS.n744 VSS.n724 5.27109
R3905 VSS.n696 VSS.n683 5.27109
R3906 VSS.n1009 VSS.n988 5.27109
R3907 VSS.n961 VSS.n960 5.27109
R3908 VSS.n906 VSS.t11 5.21007
R3909 VSS.n1829 VSS.t14 5.21007
R3910 VSS.n2457 VSS.n2456 5.0877
R3911 VSS.n2198 VSS.n2197 4.68911
R3912 VSS.n1612 VSS.t51 4.68911
R3913 VSS.n1573 VSS.n1571 4.5683
R3914 VSS.n2055 VSS.n2054 4.5683
R3915 VSS.n389 VSS.n388 4.51815
R3916 VSS.n2405 VSS.n76 4.51815
R3917 VSS.n1574 VSS.n1573 4.5005
R3918 VSS.n2054 VSS.n2053 4.5005
R3919 VSS.n2456 VSS.n73 4.26732
R3920 VSS.n2102 VSS.n519 4.19219
R3921 VSS.n1372 VSS.n1150 4.16815
R3922 VSS.n32 VSS.n3 3.81995
R3923 VSS.n318 VSS.n292 3.76521
R3924 VSS.n290 VSS.n288 3.76521
R3925 VSS.n295 VSS.n294 3.76521
R3926 VSS.n365 VSS.n363 3.76521
R3927 VSS.n378 VSS.n367 3.76521
R3928 VSS.n350 VSS.n349 3.76521
R3929 VSS.n69 VSS.n45 3.76521
R3930 VSS.n56 VSS.n50 3.76521
R3931 VSS.n28 VSS.n5 3.76521
R3932 VSS.n15 VSS.n14 3.76521
R3933 VSS.n1473 VSS.n1472 3.76521
R3934 VSS.n748 VSS.n747 3.76521
R3935 VSS.n695 VSS.n685 3.76521
R3936 VSS.n1010 VSS.n986 3.76521
R3937 VSS.n957 VSS.n948 3.76521
R3938 VSS.n1566 VSS.t79 3.6472
R3939 VSS.n1580 VSS.t13 3.6472
R3940 VSS.n1569 VSS.n1568 3.38874
R3941 VSS.n2058 VSS.n2057 3.38874
R3942 VSS.n386 VSS.n385 3.11834
R3943 VSS.n731 VSS.n729 3.09986
R3944 VSS.n711 VSS.n678 3.09986
R3945 VSS.n996 VSS.n995 3.09986
R3946 VSS.n971 VSS.n940 3.09986
R3947 VSS.n1033 VSS.n1032 3.01226
R3948 VSS.n2059 VSS.n666 3.01226
R3949 VSS VSS.n2458 2.95131
R3950 VSS.n324 VSS.n323 2.89851
R3951 VSS.n368 VSS.n347 2.89851
R3952 VSS.n51 VSS.n43 2.67025
R3953 VSS.n73 VSS.n72 2.67025
R3954 VSS.n32 VSS.n31 2.67025
R3955 VSS.n1386 VSS.t36 2.60528
R3956 VSS.n873 VSS.t19 2.60528
R3957 VSS.n1572 VSS.n519 2.5952
R3958 VSS.t85 VSS.n760 2.48621
R3959 VSS.n760 VSS.t82 2.48621
R3960 VSS.t69 VSS.n761 2.48621
R3961 VSS.n761 VSS.t85 2.48621
R3962 VSS.t52 VSS.n762 2.48621
R3963 VSS.n762 VSS.t69 2.48621
R3964 VSS.t102 VSS.n763 2.48621
R3965 VSS.n763 VSS.t52 2.48621
R3966 VSS.n712 VSS.t37 2.48621
R3967 VSS.t54 VSS.n712 2.48621
R3968 VSS.n713 VSS.t54 2.48621
R3969 VSS.n713 VSS.t75 2.48621
R3970 VSS.n716 VSS.t75 2.48621
R3971 VSS.t94 VSS.n716 2.48621
R3972 VSS.n717 VSS.t94 2.48621
R3973 VSS.t90 VSS.n717 2.48621
R3974 VSS.n764 VSS.t90 2.48621
R3975 VSS.n764 VSS.t102 2.48621
R3976 VSS.t92 VSS.n1023 2.48621
R3977 VSS.n1023 VSS.t42 2.48621
R3978 VSS.t71 VSS.n1024 2.48621
R3979 VSS.n1024 VSS.t92 2.48621
R3980 VSS.t73 VSS.n1025 2.48621
R3981 VSS.n1025 VSS.t71 2.48621
R3982 VSS.t77 VSS.n1026 2.48621
R3983 VSS.n1026 VSS.t73 2.48621
R3984 VSS.n975 VSS.t45 2.48621
R3985 VSS.t40 VSS.n975 2.48621
R3986 VSS.n976 VSS.t40 2.48621
R3987 VSS.n976 VSS.t34 2.48621
R3988 VSS.n979 VSS.t34 2.48621
R3989 VSS.t104 VSS.n979 2.48621
R3990 VSS.n980 VSS.t104 2.48621
R3991 VSS.t80 VSS.n980 2.48621
R3992 VSS.n1027 VSS.t80 2.48621
R3993 VSS.n1027 VSS.t77 2.48621
R3994 VSS.n2455 VSS.n2454 2.33344
R3995 VSS.n299 VSS.n296 2.25932
R3996 VSS.n354 VSS.n351 2.25932
R3997 VSS.n68 VSS.n47 2.25932
R3998 VSS.n18 VSS.n10 2.25932
R3999 VSS.n751 VSS.n722 2.25932
R4000 VSS.n692 VSS.n691 2.25932
R4001 VSS.n1014 VSS.n1013 2.25932
R4002 VSS.n956 VSS.n950 2.25932
R4003 VSS.n307 VSS.n74 2.25177
R4004 VSS.n385 VSS.n384 2.25177
R4005 VSS.n1580 VSS.t110 2.08433
R4006 VSS.n1667 VSS.t2 2.08433
R4007 VSS.n2458 VSS.n2457 1.74238
R4008 VSS.n429 VSS.t59 1.56337
R4009 VSS.t47 VSS.n104 1.56337
R4010 VSS.n1493 VSS.t10 1.56337
R4011 VSS.n34 VSS.n32 1.1502
R4012 VSS.n36 VSS.n34 1.1502
R4013 VSS.n38 VSS.n36 1.1502
R4014 VSS.n40 VSS.n38 1.1502
R4015 VSS.n42 VSS.n40 1.1502
R4016 VSS.n43 VSS.n42 1.1502
R4017 VSS.n73 VSS.n43 1.1502
R4018 VSS.n1382 VSS.t30 1.04241
R4019 VSS.n2456 VSS.n2455 0.805174
R4020 VSS.n2455 VSS.n74 0.7864
R4021 VSS.n759 VSS.n754 0.779912
R4022 VSS.n759 VSS.n719 0.779912
R4023 VSS.n719 VSS.n718 0.779912
R4024 VSS.n718 VSS.n671 0.779912
R4025 VSS.n688 VSS.n676 0.779912
R4026 VSS.n714 VSS.n676 0.779912
R4027 VSS.n715 VSS.n714 0.779912
R4028 VSS.n715 VSS.n670 0.779912
R4029 VSS.n765 VSS.n670 0.779912
R4030 VSS.n765 VSS.n671 0.779912
R4031 VSS.n1022 VSS.n1017 0.779912
R4032 VSS.n1022 VSS.n982 0.779912
R4033 VSS.n982 VSS.n981 0.779912
R4034 VSS.n981 VSS.n934 0.779912
R4035 VSS.n951 VSS.n939 0.779912
R4036 VSS.n977 VSS.n939 0.779912
R4037 VSS.n978 VSS.n977 0.779912
R4038 VSS.n978 VSS.n933 0.779912
R4039 VSS.n1028 VSS.n933 0.779912
R4040 VSS.n1028 VSS.n934 0.779912
R4041 VSS.n65 VSS.n64 0.753441
R4042 VSS.n20 VSS.n19 0.753441
R4043 VSS.n285 VSS.n284 0.753441
R4044 VSS.n2408 VSS.n2404 0.753441
R4045 VSS.n1471 VSS.n1470 0.753441
R4046 VSS.n1582 VSS.n1031 0.753441
R4047 VSS.n2051 VSS.n769 0.753441
R4048 VSS.n755 VSS.n668 0.701719
R4049 VSS.n756 VSS.n755 0.701719
R4050 VSS.n757 VSS.n756 0.701719
R4051 VSS.n674 VSS.n673 0.701719
R4052 VSS.n673 VSS.n672 0.701719
R4053 VSS.n672 VSS.n669 0.701719
R4054 VSS.n1018 VSS.n931 0.701719
R4055 VSS.n1019 VSS.n1018 0.701719
R4056 VSS.n1020 VSS.n1019 0.701719
R4057 VSS.n937 VSS.n936 0.701719
R4058 VSS.n936 VSS.n935 0.701719
R4059 VSS.n935 VSS.n932 0.701719
R4060 VSS.n308 VSS.n307 0.647239
R4061 VSS.n384 VSS.n383 0.647239
R4062 VSS.n1572 VSS.n0 0.633833
R4063 VSS.n385 VSS.n347 0.574311
R4064 VSS.n347 VSS.n346 0.574311
R4065 VSS.n346 VSS.n344 0.574311
R4066 VSS.n344 VSS.n342 0.574311
R4067 VSS.n342 VSS.n340 0.574311
R4068 VSS.n340 VSS.n338 0.574311
R4069 VSS.n338 VSS.n336 0.574311
R4070 VSS.n336 VSS.n334 0.574311
R4071 VSS.n334 VSS.n332 0.574311
R4072 VSS.n332 VSS.n330 0.574311
R4073 VSS.n330 VSS.n328 0.574311
R4074 VSS.n328 VSS.n326 0.574311
R4075 VSS.n326 VSS.n324 0.574311
R4076 VSS.n324 VSS.n74 0.574311
R4077 VSS.n2249 VSS.t28 0.521457
R4078 VSS.n2310 VSS.t15 0.521457
R4079 VSS.n307 VSS.n306 0.418978
R4080 VSS.n384 VSS.n361 0.418978
R4081 VSS.n758 VSS.n757 0.35111
R4082 VSS.n675 VSS.n674 0.35111
R4083 VSS.n1021 VSS.n1020 0.35111
R4084 VSS.n938 VSS.n937 0.35111
R4085 VSS.n312 VSS.n311 0.320353
R4086 VSS.n314 VSS.n312 0.320353
R4087 VSS.n314 VSS.n313 0.320353
R4088 VSS.n298 VSS.n297 0.320353
R4089 VSS.n374 VSS.n373 0.320353
R4090 VSS.n372 VSS.n369 0.320353
R4091 VSS.n373 VSS.n372 0.320353
R4092 VSS.n353 VSS.n352 0.320353
R4093 VSS.n52 VSS.n48 0.320353
R4094 VSS.n60 VSS.n48 0.320353
R4095 VSS.n61 VSS.n60 0.320353
R4096 VSS.n66 VSS.n61 0.320353
R4097 VSS.n9 VSS.n7 0.320353
R4098 VSS.n23 VSS.n7 0.320353
R4099 VSS.n24 VSS.n23 0.320353
R4100 VSS.n25 VSS.n24 0.320353
R4101 VSS VSS.n0 0.309591
R4102 VSS.n2457 VSS.n2 0.303278
R4103 VSS.n2458 VSS.n1 0.303278
R4104 VSS.n766 VSS.n765 0.272321
R4105 VSS.n1029 VSS.n1028 0.272321
R4106 VSS.n766 VSS.n668 0.261436
R4107 VSS.n766 VSS.n669 0.261436
R4108 VSS.n1029 VSS.n931 0.261436
R4109 VSS.n1029 VSS.n932 0.261436
R4110 VSS.n759 VSS.n758 0.228761
R4111 VSS.n676 VSS.n675 0.228761
R4112 VSS.n1022 VSS.n1021 0.228761
R4113 VSS.n939 VSS.n938 0.228761
R4114 VSS.n2102 VSS.n2101 0.21925
R4115 VSS.n2053 VSS.n2052 0.217762
R4116 VSS.n1575 VSS.n1574 0.217762
R4117 VSS.n2409 VSS.n75 0.204927
R4118 VSS.n387 VSS.n286 0.204927
R4119 VSS.n323 VSS.n287 0.196152
R4120 VSS.n310 VSS.n287 0.196152
R4121 VSS.n311 VSS.n310 0.196152
R4122 VSS.n301 VSS.n298 0.196152
R4123 VSS.n301 VSS.n300 0.196152
R4124 VSS.n300 VSS.n293 0.196152
R4125 VSS.n306 VSS.n293 0.196152
R4126 VSS.n317 VSS.n308 0.196152
R4127 VSS.n317 VSS.n316 0.196152
R4128 VSS.n316 VSS.n314 0.196152
R4129 VSS.n377 VSS.n368 0.196152
R4130 VSS.n377 VSS.n376 0.196152
R4131 VSS.n376 VSS.n374 0.196152
R4132 VSS.n356 VSS.n353 0.196152
R4133 VSS.n356 VSS.n355 0.196152
R4134 VSS.n355 VSS.n348 0.196152
R4135 VSS.n361 VSS.n348 0.196152
R4136 VSS.n383 VSS.n362 0.196152
R4137 VSS.n371 VSS.n362 0.196152
R4138 VSS.n372 VSS.n371 0.196152
R4139 VSS.n55 VSS.n51 0.196152
R4140 VSS.n55 VSS.n54 0.196152
R4141 VSS.n54 VSS.n52 0.196152
R4142 VSS.n72 VSS.n44 0.196152
R4143 VSS.n67 VSS.n44 0.196152
R4144 VSS.n67 VSS.n66 0.196152
R4145 VSS.n13 VSS.n3 0.196152
R4146 VSS.n13 VSS.n12 0.196152
R4147 VSS.n12 VSS.n9 0.196152
R4148 VSS.n31 VSS.n4 0.196152
R4149 VSS.n26 VSS.n4 0.196152
R4150 VSS.n26 VSS.n25 0.196152
R4151 VSS.n754 VSS.n753 0.196152
R4152 VSS.n753 VSS.n721 0.196152
R4153 VSS.n746 VSS.n721 0.196152
R4154 VSS.n746 VSS.n745 0.196152
R4155 VSS.n745 VSS.n725 0.196152
R4156 VSS.n738 VSS.n725 0.196152
R4157 VSS.n738 VSS.n737 0.196152
R4158 VSS.n737 VSS.n729 0.196152
R4159 VSS.n688 VSS.n686 0.196152
R4160 VSS.n693 VSS.n686 0.196152
R4161 VSS.n694 VSS.n693 0.196152
R4162 VSS.n694 VSS.n682 0.196152
R4163 VSS.n701 VSS.n682 0.196152
R4164 VSS.n703 VSS.n701 0.196152
R4165 VSS.n703 VSS.n702 0.196152
R4166 VSS.n702 VSS.n678 0.196152
R4167 VSS.n996 VSS.n991 0.196152
R4168 VSS.n1003 VSS.n991 0.196152
R4169 VSS.n1004 VSS.n1003 0.196152
R4170 VSS.n1004 VSS.n987 0.196152
R4171 VSS.n1011 VSS.n987 0.196152
R4172 VSS.n1012 VSS.n1011 0.196152
R4173 VSS.n1012 VSS.n983 0.196152
R4174 VSS.n1017 VSS.n983 0.196152
R4175 VSS.n971 VSS.n970 0.196152
R4176 VSS.n970 VSS.n943 0.196152
R4177 VSS.n963 VSS.n943 0.196152
R4178 VSS.n963 VSS.n962 0.196152
R4179 VSS.n962 VSS.n947 0.196152
R4180 VSS.n955 VSS.n947 0.196152
R4181 VSS.n955 VSS.n954 0.196152
R4182 VSS.n954 VSS.n951 0.196152
R4183 VSS.n1571 VSS.n1570 0.193208
R4184 VSS.n2056 VSS.n2055 0.193208
R4185 VSS.n1793 VSS.n0 0.172159
R4186 VSS.n767 VSS.n766 0.114136
R4187 VSS.n1030 VSS.n1029 0.114136
R4188 VSS.n2454 VSS.n75 0.104667
R4189 VSS.n387 VSS.n386 0.104667
R4190 VSS.n1571 VSS.n1030 0.048119
R4191 VSS.n1574 VSS.n1030 0.048119
R4192 VSS.n2055 VSS.n767 0.048119
R4193 VSS.n2053 VSS.n767 0.048119
R4194 a_2479_7336.n1 a_2479_7336.t31 260.486
R4195 a_2479_7336.n11 a_2479_7336.t19 260.486
R4196 a_2479_7336.n9 a_2479_7336.t34 260.111
R4197 a_2479_7336.n8 a_2479_7336.t21 260.111
R4198 a_2479_7336.n7 a_2479_7336.t29 260.111
R4199 a_2479_7336.n6 a_2479_7336.t18 260.111
R4200 a_2479_7336.n5 a_2479_7336.t33 260.111
R4201 a_2479_7336.n4 a_2479_7336.t27 260.111
R4202 a_2479_7336.n2 a_2479_7336.t24 260.111
R4203 a_2479_7336.n1 a_2479_7336.t22 260.111
R4204 a_2479_7336.n11 a_2479_7336.t28 260.111
R4205 a_2479_7336.n12 a_2479_7336.t35 260.111
R4206 a_2479_7336.n14 a_2479_7336.t32 260.111
R4207 a_2479_7336.n15 a_2479_7336.t26 260.111
R4208 a_2479_7336.n16 a_2479_7336.t23 260.111
R4209 a_2479_7336.n17 a_2479_7336.t20 260.111
R4210 a_2479_7336.n18 a_2479_7336.t30 260.111
R4211 a_2479_7336.n19 a_2479_7336.t25 260.111
R4212 a_2479_7336.n3 a_2479_7336.n0 203.843
R4213 a_2479_7336.n13 a_2479_7336.n10 203.843
R4214 a_2479_7336.n81 a_2479_7336.n63 185
R4215 a_2479_7336.n81 a_2479_7336.n62 185
R4216 a_2479_7336.n81 a_2479_7336.n61 185
R4217 a_2479_7336.n81 a_2479_7336.n60 185
R4218 a_2479_7336.n81 a_2479_7336.n59 185
R4219 a_2479_7336.n81 a_2479_7336.n58 185
R4220 a_2479_7336.n81 a_2479_7336.n57 185
R4221 a_2479_7336.n50 a_2479_7336.n32 185
R4222 a_2479_7336.n50 a_2479_7336.n31 185
R4223 a_2479_7336.n50 a_2479_7336.n30 185
R4224 a_2479_7336.n50 a_2479_7336.n29 185
R4225 a_2479_7336.n50 a_2479_7336.n28 185
R4226 a_2479_7336.n50 a_2479_7336.n27 185
R4227 a_2479_7336.n50 a_2479_7336.n26 185
R4228 a_2479_7336.n65 a_2479_7336.t4 130.75
R4229 a_2479_7336.n34 a_2479_7336.t7 130.75
R4230 a_2479_7336.n65 a_2479_7336.t6 91.3557
R4231 a_2479_7336.n34 a_2479_7336.t8 91.3557
R4232 a_2479_7336.n82 a_2479_7336.n81 86.5152
R4233 a_2479_7336.n51 a_2479_7336.n50 86.5152
R4234 a_2479_7336.n80 a_2479_7336.n64 30.3012
R4235 a_2479_7336.n49 a_2479_7336.n33 30.3012
R4236 a_2479_7336.n0 a_2479_7336.t13 28.5655
R4237 a_2479_7336.n0 a_2479_7336.t14 28.5655
R4238 a_2479_7336.n10 a_2479_7336.t15 28.5655
R4239 a_2479_7336.n10 a_2479_7336.t3 28.5655
R4240 a_2479_7336.n57 a_2479_7336.n56 24.8476
R4241 a_2479_7336.n26 a_2479_7336.n25 24.8476
R4242 a_2479_7336.n66 a_2479_7336.n58 23.3417
R4243 a_2479_7336.n35 a_2479_7336.n27 23.3417
R4244 a_2479_7336.n83 a_2479_7336.n82 22.0256
R4245 a_2479_7336.n52 a_2479_7336.n51 22.0256
R4246 a_2479_7336.n68 a_2479_7336.n59 21.8358
R4247 a_2479_7336.n37 a_2479_7336.n28 21.8358
R4248 a_2479_7336.n70 a_2479_7336.n60 20.3299
R4249 a_2479_7336.n39 a_2479_7336.n29 20.3299
R4250 a_2479_7336.n72 a_2479_7336.n61 18.824
R4251 a_2479_7336.n41 a_2479_7336.n30 18.824
R4252 a_2479_7336.n74 a_2479_7336.n62 17.3181
R4253 a_2479_7336.n43 a_2479_7336.n31 17.3181
R4254 a_2479_7336.n81 a_2479_7336.n80 16.3559
R4255 a_2479_7336.n50 a_2479_7336.n49 16.3559
R4256 a_2479_7336.n76 a_2479_7336.n63 15.8123
R4257 a_2479_7336.n45 a_2479_7336.n32 15.8123
R4258 a_2479_7336.n86 a_2479_7336.n85 14.6053
R4259 a_2479_7336.n23 a_2479_7336.n22 14.6052
R4260 a_2479_7336.n54 a_2479_7336.n53 14.377
R4261 a_2479_7336.n82 a_2479_7336.n56 12.7256
R4262 a_2479_7336.n51 a_2479_7336.n25 12.7256
R4263 a_2479_7336.n20 a_2479_7336.t17 12.5928
R4264 a_2479_7336.n85 a_2479_7336.n84 11.5586
R4265 a_2479_7336.n64 a_2479_7336.n63 11.2946
R4266 a_2479_7336.n33 a_2479_7336.n32 11.2946
R4267 a_2479_7336.n76 a_2479_7336.n62 9.78874
R4268 a_2479_7336.n45 a_2479_7336.n31 9.78874
R4269 a_2479_7336.n56 a_2479_7336.n55 9.3005
R4270 a_2479_7336.n67 a_2479_7336.n66 9.3005
R4271 a_2479_7336.n69 a_2479_7336.n68 9.3005
R4272 a_2479_7336.n71 a_2479_7336.n70 9.3005
R4273 a_2479_7336.n73 a_2479_7336.n72 9.3005
R4274 a_2479_7336.n75 a_2479_7336.n74 9.3005
R4275 a_2479_7336.n77 a_2479_7336.n76 9.3005
R4276 a_2479_7336.n78 a_2479_7336.n64 9.3005
R4277 a_2479_7336.n25 a_2479_7336.n24 9.3005
R4278 a_2479_7336.n36 a_2479_7336.n35 9.3005
R4279 a_2479_7336.n38 a_2479_7336.n37 9.3005
R4280 a_2479_7336.n40 a_2479_7336.n39 9.3005
R4281 a_2479_7336.n42 a_2479_7336.n41 9.3005
R4282 a_2479_7336.n44 a_2479_7336.n43 9.3005
R4283 a_2479_7336.n46 a_2479_7336.n45 9.3005
R4284 a_2479_7336.n47 a_2479_7336.n33 9.3005
R4285 a_2479_7336.n74 a_2479_7336.n61 8.28285
R4286 a_2479_7336.n43 a_2479_7336.n30 8.28285
R4287 a_2479_7336.n23 a_2479_7336.n21 8.22405
R4288 a_2479_7336.n72 a_2479_7336.n60 6.77697
R4289 a_2479_7336.n41 a_2479_7336.n29 6.77697
R4290 a_2479_7336.n54 a_2479_7336.n52 6.19091
R4291 a_2479_7336.n70 a_2479_7336.n59 5.27109
R4292 a_2479_7336.n39 a_2479_7336.n28 5.27109
R4293 a_2479_7336.n21 a_2479_7336.n20 4.66982
R4294 a_2479_7336.n68 a_2479_7336.n58 3.76521
R4295 a_2479_7336.n37 a_2479_7336.n27 3.76521
R4296 a_2479_7336.n84 a_2479_7336.n83 3.31388
R4297 a_2479_7336.n85 a_2479_7336.n23 2.87753
R4298 a_2479_7336.n22 a_2479_7336.t2 2.48621
R4299 a_2479_7336.n22 a_2479_7336.t1 2.48621
R4300 a_2479_7336.n81 a_2479_7336.t10 2.48621
R4301 a_2479_7336.n81 a_2479_7336.t5 2.48621
R4302 a_2479_7336.n50 a_2479_7336.t8 2.48621
R4303 a_2479_7336.n50 a_2479_7336.t12 2.48621
R4304 a_2479_7336.n53 a_2479_7336.t9 2.48621
R4305 a_2479_7336.n53 a_2479_7336.t16 2.48621
R4306 a_2479_7336.n86 a_2479_7336.t11 2.48621
R4307 a_2479_7336.t0 a_2479_7336.n86 2.48621
R4308 a_2479_7336.n80 a_2479_7336.n79 2.36936
R4309 a_2479_7336.n49 a_2479_7336.n48 2.36936
R4310 a_2479_7336.n84 a_2479_7336.n54 2.30287
R4311 a_2479_7336.n66 a_2479_7336.n57 2.25932
R4312 a_2479_7336.n35 a_2479_7336.n26 2.25932
R4313 a_2479_7336.n20 a_2479_7336.n19 1.41083
R4314 a_2479_7336.n21 a_2479_7336.n9 1.3088
R4315 a_2479_7336.n2 a_2479_7336.n1 0.3755
R4316 a_2479_7336.n5 a_2479_7336.n4 0.3755
R4317 a_2479_7336.n6 a_2479_7336.n5 0.3755
R4318 a_2479_7336.n7 a_2479_7336.n6 0.3755
R4319 a_2479_7336.n8 a_2479_7336.n7 0.3755
R4320 a_2479_7336.n9 a_2479_7336.n8 0.3755
R4321 a_2479_7336.n19 a_2479_7336.n18 0.3755
R4322 a_2479_7336.n18 a_2479_7336.n17 0.3755
R4323 a_2479_7336.n17 a_2479_7336.n16 0.3755
R4324 a_2479_7336.n16 a_2479_7336.n15 0.3755
R4325 a_2479_7336.n15 a_2479_7336.n14 0.3755
R4326 a_2479_7336.n12 a_2479_7336.n11 0.3755
R4327 a_2479_7336.n79 a_2479_7336.n65 0.320353
R4328 a_2479_7336.n48 a_2479_7336.n34 0.320353
R4329 a_2479_7336.n79 a_2479_7336.n78 0.196152
R4330 a_2479_7336.n78 a_2479_7336.n77 0.196152
R4331 a_2479_7336.n77 a_2479_7336.n75 0.196152
R4332 a_2479_7336.n75 a_2479_7336.n73 0.196152
R4333 a_2479_7336.n73 a_2479_7336.n71 0.196152
R4334 a_2479_7336.n71 a_2479_7336.n69 0.196152
R4335 a_2479_7336.n69 a_2479_7336.n67 0.196152
R4336 a_2479_7336.n67 a_2479_7336.n55 0.196152
R4337 a_2479_7336.n83 a_2479_7336.n55 0.196152
R4338 a_2479_7336.n48 a_2479_7336.n47 0.196152
R4339 a_2479_7336.n47 a_2479_7336.n46 0.196152
R4340 a_2479_7336.n46 a_2479_7336.n44 0.196152
R4341 a_2479_7336.n44 a_2479_7336.n42 0.196152
R4342 a_2479_7336.n42 a_2479_7336.n40 0.196152
R4343 a_2479_7336.n40 a_2479_7336.n38 0.196152
R4344 a_2479_7336.n38 a_2479_7336.n36 0.196152
R4345 a_2479_7336.n36 a_2479_7336.n24 0.196152
R4346 a_2479_7336.n52 a_2479_7336.n24 0.196152
R4347 a_2479_7336.n3 a_2479_7336.n2 0.188
R4348 a_2479_7336.n4 a_2479_7336.n3 0.188
R4349 a_2479_7336.n14 a_2479_7336.n13 0.188
R4350 a_2479_7336.n13 a_2479_7336.n12 0.188
R4351 VOUT.n13 VOUT.t26 260.298
R4352 VOUT.t22 VOUT.n13 260.298
R4353 VOUT.t26 VOUT.n8 260.298
R4354 VOUT.n50 VOUT.t24 260.298
R4355 VOUT.t20 VOUT.n50 260.298
R4356 VOUT.n51 VOUT.t20 260.298
R4357 VOUT.n14 VOUT.t22 260.111
R4358 VOUT.t24 VOUT.n48 260.111
R4359 VOUT.n12 VOUT.t28 232.03
R4360 VOUT.t21 VOUT.n49 232.03
R4361 VOUT.n2 VOUT.n0 206.708
R4362 VOUT.n6 VOUT.n5 206.094
R4363 VOUT.n4 VOUT.n3 206.094
R4364 VOUT.n2 VOUT.n1 206.094
R4365 VOUT.n64 VOUT.n63 206.094
R4366 VOUT.n62 VOUT.n61 206.094
R4367 VOUT.n60 VOUT.n59 206.094
R4368 VOUT.n58 VOUT.n57 206.094
R4369 VOUT.n11 VOUT.n10 203.03
R4370 VOUT.n9 VOUT.n7 203.03
R4371 VOUT.n55 VOUT.n54 203.03
R4372 VOUT.n53 VOUT.n52 203.03
R4373 VOUT.n43 VOUT.n42 185
R4374 VOUT.n43 VOUT.n25 185
R4375 VOUT.n43 VOUT.n24 185
R4376 VOUT.n43 VOUT.n23 185
R4377 VOUT.n43 VOUT.n22 185
R4378 VOUT.n43 VOUT.n21 185
R4379 VOUT.n43 VOUT.n20 185
R4380 VOUT.n26 VOUT.t29 130.75
R4381 VOUT.n26 VOUT.t31 91.3557
R4382 VOUT.n44 VOUT.n43 86.5152
R4383 VOUT.n28 VOUT.n19 30.3012
R4384 VOUT.n10 VOUT.t23 28.5655
R4385 VOUT.n10 VOUT.t27 28.5655
R4386 VOUT.n9 VOUT.t12 28.5655
R4387 VOUT.t23 VOUT.n9 28.5655
R4388 VOUT.n5 VOUT.t10 28.5655
R4389 VOUT.n5 VOUT.t5 28.5655
R4390 VOUT.n3 VOUT.t13 28.5655
R4391 VOUT.n3 VOUT.t7 28.5655
R4392 VOUT.n1 VOUT.t14 28.5655
R4393 VOUT.n1 VOUT.t1 28.5655
R4394 VOUT.n0 VOUT.t3 28.5655
R4395 VOUT.n0 VOUT.t8 28.5655
R4396 VOUT.n54 VOUT.t25 28.5655
R4397 VOUT.n54 VOUT.t18 28.5655
R4398 VOUT.n53 VOUT.t21 28.5655
R4399 VOUT.t25 VOUT.n53 28.5655
R4400 VOUT.n63 VOUT.t6 28.5655
R4401 VOUT.n63 VOUT.t17 28.5655
R4402 VOUT.n61 VOUT.t16 28.5655
R4403 VOUT.n61 VOUT.t9 28.5655
R4404 VOUT.n59 VOUT.t4 28.5655
R4405 VOUT.n59 VOUT.t15 28.5655
R4406 VOUT.n57 VOUT.t2 28.5655
R4407 VOUT.n57 VOUT.t11 28.5655
R4408 VOUT.n42 VOUT.n18 24.8476
R4409 VOUT.n41 VOUT.n25 23.3417
R4410 VOUT.n45 VOUT.n44 22.0256
R4411 VOUT.n38 VOUT.n24 21.8358
R4412 VOUT.n36 VOUT.n23 20.3299
R4413 VOUT.n46 VOUT.n45 19.0885
R4414 VOUT.n34 VOUT.n22 18.824
R4415 VOUT.n32 VOUT.n21 17.3181
R4416 VOUT.n43 VOUT.n19 16.3559
R4417 VOUT.n30 VOUT.n20 15.8123
R4418 VOUT.n44 VOUT.n18 12.7256
R4419 VOUT.n28 VOUT.n20 11.2946
R4420 VOUT.n30 VOUT.n21 9.78874
R4421 VOUT.n18 VOUT.n17 9.3005
R4422 VOUT.n41 VOUT.n40 9.3005
R4423 VOUT.n39 VOUT.n38 9.3005
R4424 VOUT.n37 VOUT.n36 9.3005
R4425 VOUT.n35 VOUT.n34 9.3005
R4426 VOUT.n33 VOUT.n32 9.3005
R4427 VOUT.n31 VOUT.n30 9.3005
R4428 VOUT.n29 VOUT.n28 9.3005
R4429 VOUT.n32 VOUT.n22 8.28285
R4430 VOUT.n34 VOUT.n23 6.77697
R4431 VOUT.n36 VOUT.n24 5.27109
R4432 VOUT.n47 VOUT.t19 3.9533
R4433 VOUT.n38 VOUT.n25 3.76521
R4434 VOUT.n66 VOUT.n46 3.29996
R4435 VOUT.n58 VOUT.n56 3.23261
R4436 VOUT.n16 VOUT.n15 2.55612
R4437 VOUT.n43 VOUT.t0 2.48621
R4438 VOUT.n43 VOUT.t30 2.48621
R4439 VOUT VOUT.n16 2.47337
R4440 VOUT.n27 VOUT.n19 2.36936
R4441 VOUT.n42 VOUT.n41 2.25932
R4442 VOUT.n65 VOUT.n64 2.12962
R4443 VOUT.n66 VOUT.n65 1.09816
R4444 VOUT.n4 VOUT.n2 0.61449
R4445 VOUT.n6 VOUT.n4 0.61449
R4446 VOUT.n16 VOUT.n6 0.61449
R4447 VOUT.n60 VOUT.n58 0.61449
R4448 VOUT.n62 VOUT.n60 0.61449
R4449 VOUT.n64 VOUT.n62 0.61449
R4450 VOUT VOUT.n66 0.521984
R4451 VOUT.n56 VOUT.n55 0.446229
R4452 VOUT.n55 VOUT.n49 0.43664
R4453 VOUT.n12 VOUT.n7 0.436638
R4454 VOUT.n15 VOUT.n7 0.38373
R4455 VOUT.n11 VOUT.n8 0.38373
R4456 VOUT.n52 VOUT.n51 0.383729
R4457 VOUT.n27 VOUT.n26 0.320353
R4458 VOUT.n13 VOUT.n12 0.285826
R4459 VOUT.n50 VOUT.n49 0.285826
R4460 VOUT.n47 VOUT.n46 0.220947
R4461 VOUT.n45 VOUT.n17 0.196152
R4462 VOUT.n40 VOUT.n17 0.196152
R4463 VOUT.n40 VOUT.n39 0.196152
R4464 VOUT.n39 VOUT.n37 0.196152
R4465 VOUT.n37 VOUT.n35 0.196152
R4466 VOUT.n35 VOUT.n33 0.196152
R4467 VOUT.n33 VOUT.n31 0.196152
R4468 VOUT.n31 VOUT.n29 0.196152
R4469 VOUT.n29 VOUT.n27 0.196152
R4470 VOUT.n15 VOUT.n14 0.188
R4471 VOUT.n14 VOUT.n8 0.188
R4472 VOUT.n51 VOUT.n48 0.188
R4473 VOUT.n56 VOUT.n48 0.1255
R4474 VOUT.n52 VOUT.n49 0.0984044
R4475 VOUT.n12 VOUT.n11 0.0984028
R4476 VOUT.n65 VOUT.n47 0.0649934
R4477 VDD.n297 VDD.n68 723.529
R4478 VDD.n73 VDD.n65 723.529
R4479 VDD.n136 VDD.n112 723.529
R4480 VDD.n180 VDD.n114 723.529
R4481 VDD.n257 VDD.n256 515.294
R4482 VDD.n55 VDD.n51 275.295
R4483 VDD.n147 VDD.n131 275.295
R4484 VDD.n34 VDD.t49 260.486
R4485 VDD.n20 VDD.t24 260.486
R4486 VDD.n330 VDD.t13 260.486
R4487 VDD.n315 VDD.t33 260.486
R4488 VDD.t6 VDD.n38 260.298
R4489 VDD.n36 VDD.t27 260.298
R4490 VDD.n39 VDD.t6 260.298
R4491 VDD.t46 VDD.n19 260.298
R4492 VDD.n17 VDD.t35 260.298
R4493 VDD.n13 VDD.t35 260.298
R4494 VDD.t19 VDD.n327 260.298
R4495 VDD.t37 VDD.n329 260.298
R4496 VDD.n334 VDD.t19 260.298
R4497 VDD.n312 VDD.t44 260.298
R4498 VDD.t44 VDD.n309 260.298
R4499 VDD.n316 VDD.t51 260.298
R4500 VDD.n1 VDD.t16 260.199
R4501 VDD.n352 VDD.t39 260.199
R4502 VDD.t30 VDD.n32 260.111
R4503 VDD.n37 VDD.t30 260.111
R4504 VDD.t27 VDD.n34 260.111
R4505 VDD.n20 VDD.t46 260.111
R4506 VDD.t10 VDD.n12 260.111
R4507 VDD.n18 VDD.t10 260.111
R4508 VDD.n333 VDD.t42 260.111
R4509 VDD.t42 VDD.n332 260.111
R4510 VDD.n330 VDD.t37 260.111
R4511 VDD.t51 VDD.n315 260.111
R4512 VDD.n314 VDD.t22 260.111
R4513 VDD.t22 VDD.n313 260.111
R4514 VDD.n67 VDD.n66 240
R4515 VDD.n292 VDD.n66 240
R4516 VDD.n290 VDD.n289 240
R4517 VDD.n301 VDD.n50 240
R4518 VDD.n253 VDD.n252 240
R4519 VDD.n261 VDD.n260 240
R4520 VDD.n265 VDD.n264 240
R4521 VDD.n269 VDD.n268 240
R4522 VDD.n273 VDD.n272 240
R4523 VDD.n277 VDD.n276 240
R4524 VDD.n279 VDD.n65 240
R4525 VDD.n186 VDD.n112 240
R4526 VDD.n186 VDD.n110 240
R4527 VDD.n190 VDD.n110 240
R4528 VDD.n190 VDD.n105 240
R4529 VDD.n199 VDD.n105 240
R4530 VDD.n199 VDD.n103 240
R4531 VDD.n203 VDD.n103 240
R4532 VDD.n203 VDD.n98 240
R4533 VDD.n212 VDD.n98 240
R4534 VDD.n212 VDD.n96 240
R4535 VDD.n216 VDD.n96 240
R4536 VDD.n216 VDD.n91 240
R4537 VDD.n224 VDD.n91 240
R4538 VDD.n224 VDD.n89 240
R4539 VDD.n228 VDD.n89 240
R4540 VDD.n228 VDD.n83 240
R4541 VDD.n236 VDD.n83 240
R4542 VDD.n236 VDD.n81 240
R4543 VDD.n240 VDD.n81 240
R4544 VDD.n240 VDD.n75 240
R4545 VDD.n248 VDD.n75 240
R4546 VDD.n248 VDD.n72 240
R4547 VDD.n284 VDD.n72 240
R4548 VDD.n284 VDD.n73 240
R4549 VDD.n178 VDD.n177 240
R4550 VDD.n175 VDD.n119 240
R4551 VDD.n171 VDD.n170 240
R4552 VDD.n168 VDD.n122 240
R4553 VDD.n164 VDD.n163 240
R4554 VDD.n161 VDD.n125 240
R4555 VDD.n157 VDD.n156 240
R4556 VDD.n154 VDD.n128 240
R4557 VDD.n150 VDD.n149 240
R4558 VDD.n143 VDD.n142 240
R4559 VDD.n140 VDD.n134 240
R4560 VDD.n184 VDD.n114 240
R4561 VDD.n184 VDD.n109 240
R4562 VDD.n193 VDD.n109 240
R4563 VDD.n193 VDD.n107 240
R4564 VDD.n197 VDD.n107 240
R4565 VDD.n197 VDD.n102 240
R4566 VDD.n206 VDD.n102 240
R4567 VDD.n206 VDD.n100 240
R4568 VDD.n210 VDD.n100 240
R4569 VDD.n210 VDD.n95 240
R4570 VDD.n218 VDD.n95 240
R4571 VDD.n218 VDD.n93 240
R4572 VDD.n222 VDD.n93 240
R4573 VDD.n222 VDD.n87 240
R4574 VDD.n230 VDD.n87 240
R4575 VDD.n230 VDD.n85 240
R4576 VDD.n234 VDD.n85 240
R4577 VDD.n234 VDD.n79 240
R4578 VDD.n242 VDD.n79 240
R4579 VDD.n242 VDD.n77 240
R4580 VDD.n246 VDD.n77 240
R4581 VDD.n246 VDD.n70 240
R4582 VDD.n286 VDD.n70 240
R4583 VDD.n286 VDD.n68 240
R4584 VDD.n31 VDD.t9 232.03
R4585 VDD.n16 VDD.t36 232.03
R4586 VDD.n335 VDD.t21 232.03
R4587 VDD.t45 VDD.n308 232.03
R4588 VDD.n351 VDD.t41 231.758
R4589 VDD.n345 VDD.n343 206.48
R4590 VDD.n324 VDD.n323 205.865
R4591 VDD.n349 VDD.n348 205.865
R4592 VDD.n347 VDD.n346 205.865
R4593 VDD.n345 VDD.n344 205.865
R4594 VDD.n9 VDD.n8 205.865
R4595 VDD.n7 VDD.n6 205.865
R4596 VDD.n5 VDD.n4 205.865
R4597 VDD.n3 VDD.n2 205.865
R4598 VDD.n28 VDD.n27 205.865
R4599 VDD.n351 VDD.n350 203.143
R4600 VDD.n45 VDD.n44 203.127
R4601 VDD.n26 VDD.n25 203.127
R4602 VDD.n341 VDD.n340 203.127
R4603 VDD.n322 VDD.n321 203.127
R4604 VDD.n43 VDD.n29 203.126
R4605 VDD.n24 VDD.n10 203.126
R4606 VDD.n339 VDD.n325 203.126
R4607 VDD.n320 VDD.n306 203.126
R4608 VDD.n42 VDD.n30 203.03
R4609 VDD.n41 VDD.n40 203.03
R4610 VDD.n23 VDD.n22 203.03
R4611 VDD.n15 VDD.n14 203.03
R4612 VDD.n338 VDD.n326 203.03
R4613 VDD.n337 VDD.n336 203.03
R4614 VDD.n319 VDD.n318 203.03
R4615 VDD.n311 VDD.n310 203.03
R4616 VDD.n182 VDD.n114 185
R4617 VDD.n116 VDD.n114 185
R4618 VDD.n184 VDD.n183 185
R4619 VDD.n185 VDD.n184 185
R4620 VDD.n109 VDD.n108 185
R4621 VDD.n113 VDD.n109 185
R4622 VDD.n194 VDD.n193 185
R4623 VDD.n193 VDD.n192 185
R4624 VDD.n195 VDD.n107 185
R4625 VDD.n191 VDD.n107 185
R4626 VDD.n197 VDD.n196 185
R4627 VDD.n198 VDD.n197 185
R4628 VDD.n102 VDD.n101 185
R4629 VDD.n106 VDD.n102 185
R4630 VDD.n207 VDD.n206 185
R4631 VDD.n206 VDD.n205 185
R4632 VDD.n208 VDD.n100 185
R4633 VDD.n204 VDD.n100 185
R4634 VDD.n210 VDD.n209 185
R4635 VDD.n211 VDD.n210 185
R4636 VDD.n95 VDD.n94 185
R4637 VDD.n99 VDD.n95 185
R4638 VDD.n219 VDD.n218 185
R4639 VDD.n218 VDD.n217 185
R4640 VDD.n220 VDD.n93 185
R4641 VDD.n93 VDD.n92 185
R4642 VDD.n222 VDD.n221 185
R4643 VDD.n223 VDD.n222 185
R4644 VDD.n87 VDD.n86 185
R4645 VDD.n88 VDD.n87 185
R4646 VDD.n231 VDD.n230 185
R4647 VDD.n230 VDD.n229 185
R4648 VDD.n232 VDD.n85 185
R4649 VDD.n85 VDD.n84 185
R4650 VDD.n234 VDD.n233 185
R4651 VDD.n235 VDD.n234 185
R4652 VDD.n79 VDD.n78 185
R4653 VDD.n80 VDD.n79 185
R4654 VDD.n243 VDD.n242 185
R4655 VDD.n242 VDD.n241 185
R4656 VDD.n244 VDD.n77 185
R4657 VDD.n77 VDD.n76 185
R4658 VDD.n246 VDD.n245 185
R4659 VDD.n247 VDD.n246 185
R4660 VDD.n70 VDD.n69 185
R4661 VDD.n71 VDD.n70 185
R4662 VDD.n287 VDD.n286 185
R4663 VDD.n286 VDD.n285 185
R4664 VDD.n288 VDD.n68 185
R4665 VDD.n68 VDD.n52 185
R4666 VDD.n137 VDD.n136 185
R4667 VDD.n138 VDD.n134 185
R4668 VDD.n140 VDD.n139 185
R4669 VDD.n142 VDD.n132 185
R4670 VDD.n144 VDD.n143 185
R4671 VDD.n145 VDD.n131 185
R4672 VDD.n147 VDD.n146 185
R4673 VDD.n149 VDD.n129 185
R4674 VDD.n151 VDD.n150 185
R4675 VDD.n152 VDD.n128 185
R4676 VDD.n154 VDD.n153 185
R4677 VDD.n156 VDD.n126 185
R4678 VDD.n158 VDD.n157 185
R4679 VDD.n159 VDD.n125 185
R4680 VDD.n161 VDD.n160 185
R4681 VDD.n163 VDD.n123 185
R4682 VDD.n165 VDD.n164 185
R4683 VDD.n166 VDD.n122 185
R4684 VDD.n168 VDD.n167 185
R4685 VDD.n170 VDD.n120 185
R4686 VDD.n172 VDD.n171 185
R4687 VDD.n173 VDD.n119 185
R4688 VDD.n175 VDD.n174 185
R4689 VDD.n177 VDD.n118 185
R4690 VDD.n178 VDD.n115 185
R4691 VDD.n181 VDD.n180 185
R4692 VDD.n282 VDD.n73 185
R4693 VDD.n73 VDD.n52 185
R4694 VDD.n284 VDD.n283 185
R4695 VDD.n285 VDD.n284 185
R4696 VDD.n250 VDD.n72 185
R4697 VDD.n72 VDD.n71 185
R4698 VDD.n249 VDD.n248 185
R4699 VDD.n248 VDD.n247 185
R4700 VDD.n75 VDD.n74 185
R4701 VDD.n76 VDD.n75 185
R4702 VDD.n240 VDD.n239 185
R4703 VDD.n241 VDD.n240 185
R4704 VDD.n238 VDD.n81 185
R4705 VDD.n81 VDD.n80 185
R4706 VDD.n237 VDD.n236 185
R4707 VDD.n236 VDD.n235 185
R4708 VDD.n83 VDD.n82 185
R4709 VDD.n84 VDD.n83 185
R4710 VDD.n228 VDD.n227 185
R4711 VDD.n229 VDD.n228 185
R4712 VDD.n226 VDD.n89 185
R4713 VDD.n89 VDD.n88 185
R4714 VDD.n225 VDD.n224 185
R4715 VDD.n224 VDD.n223 185
R4716 VDD.n91 VDD.n90 185
R4717 VDD.n92 VDD.n91 185
R4718 VDD.n216 VDD.n215 185
R4719 VDD.n217 VDD.n216 185
R4720 VDD.n214 VDD.n96 185
R4721 VDD.n99 VDD.n96 185
R4722 VDD.n213 VDD.n212 185
R4723 VDD.n212 VDD.n211 185
R4724 VDD.n98 VDD.n97 185
R4725 VDD.n204 VDD.n98 185
R4726 VDD.n203 VDD.n202 185
R4727 VDD.n205 VDD.n203 185
R4728 VDD.n201 VDD.n103 185
R4729 VDD.n106 VDD.n103 185
R4730 VDD.n200 VDD.n199 185
R4731 VDD.n199 VDD.n198 185
R4732 VDD.n105 VDD.n104 185
R4733 VDD.n191 VDD.n105 185
R4734 VDD.n190 VDD.n189 185
R4735 VDD.n192 VDD.n190 185
R4736 VDD.n188 VDD.n110 185
R4737 VDD.n113 VDD.n110 185
R4738 VDD.n187 VDD.n186 185
R4739 VDD.n186 VDD.n185 185
R4740 VDD.n112 VDD.n111 185
R4741 VDD.n116 VDD.n112 185
R4742 VDD.n297 VDD.n296 185
R4743 VDD.n295 VDD.n67 185
R4744 VDD.n294 VDD.n66 185
R4745 VDD.n299 VDD.n66 185
R4746 VDD.n293 VDD.n292 185
R4747 VDD.n291 VDD.n290 185
R4748 VDD.n289 VDD.n47 185
R4749 VDD.n55 VDD.n54 185
R4750 VDD.n51 VDD.n48 185
R4751 VDD.n302 VDD.n301 185
R4752 VDD.n50 VDD.n49 185
R4753 VDD.n252 VDD.n251 185
R4754 VDD.n254 VDD.n253 185
R4755 VDD.n256 VDD.n255 185
R4756 VDD.n258 VDD.n257 185
R4757 VDD.n260 VDD.n259 185
R4758 VDD.n262 VDD.n261 185
R4759 VDD.n264 VDD.n263 185
R4760 VDD.n266 VDD.n265 185
R4761 VDD.n268 VDD.n267 185
R4762 VDD.n270 VDD.n269 185
R4763 VDD.n272 VDD.n271 185
R4764 VDD.n274 VDD.n273 185
R4765 VDD.n276 VDD.n275 185
R4766 VDD.n278 VDD.n277 185
R4767 VDD.n280 VDD.n279 185
R4768 VDD.n281 VDD.n65 185
R4769 VDD.n299 VDD.n65 185
R4770 VDD.n157 VDD.n127 107.683
R4771 VDD.n127 VDD.n125 107.683
R4772 VDD.n1 VDD.n0 101.662
R4773 VDD.n269 VDD.n62 78.9253
R4774 VDD.n169 VDD.n168 78.9253
R4775 VDD.n170 VDD.n169 78.9253
R4776 VDD.n272 VDD.n62 78.9253
R4777 VDD.n182 VDD.n181 77.177
R4778 VDD.n296 VDD.n288 77.177
R4779 VDD.n137 VDD.n111 77.177
R4780 VDD.n282 VDD.n281 77.177
R4781 VDD.n298 VDD.n297 72.7879
R4782 VDD.n292 VDD.n53 72.7879
R4783 VDD.n289 VDD.n56 72.7879
R4784 VDD.n300 VDD.n51 72.7879
R4785 VDD.n57 VDD.n50 72.7879
R4786 VDD.n253 VDD.n58 72.7879
R4787 VDD.n257 VDD.n59 72.7879
R4788 VDD.n261 VDD.n60 72.7879
R4789 VDD.n265 VDD.n61 72.7879
R4790 VDD.n273 VDD.n63 72.7879
R4791 VDD.n277 VDD.n64 72.7879
R4792 VDD.n179 VDD.n178 72.7879
R4793 VDD.n176 VDD.n175 72.7879
R4794 VDD.n171 VDD.n121 72.7879
R4795 VDD.n164 VDD.n124 72.7879
R4796 VDD.n162 VDD.n161 72.7879
R4797 VDD.n155 VDD.n154 72.7879
R4798 VDD.n150 VDD.n130 72.7879
R4799 VDD.n148 VDD.n147 72.7879
R4800 VDD.n143 VDD.n133 72.7879
R4801 VDD.n141 VDD.n140 72.7879
R4802 VDD.n136 VDD.n135 72.7879
R4803 VDD.n135 VDD.n134 72.7879
R4804 VDD.n142 VDD.n141 72.7879
R4805 VDD.n133 VDD.n131 72.7879
R4806 VDD.n149 VDD.n148 72.7879
R4807 VDD.n130 VDD.n128 72.7879
R4808 VDD.n156 VDD.n155 72.7879
R4809 VDD.n163 VDD.n162 72.7879
R4810 VDD.n124 VDD.n122 72.7879
R4811 VDD.n121 VDD.n119 72.7879
R4812 VDD.n177 VDD.n176 72.7879
R4813 VDD.n180 VDD.n179 72.7879
R4814 VDD.n298 VDD.n67 72.7879
R4815 VDD.n290 VDD.n53 72.7879
R4816 VDD.n56 VDD.n55 72.7879
R4817 VDD.n301 VDD.n300 72.7879
R4818 VDD.n252 VDD.n57 72.7879
R4819 VDD.n256 VDD.n58 72.7879
R4820 VDD.n260 VDD.n59 72.7879
R4821 VDD.n264 VDD.n60 72.7879
R4822 VDD.n268 VDD.n61 72.7879
R4823 VDD.n276 VDD.n63 72.7879
R4824 VDD.n279 VDD.n64 72.7879
R4825 VDD.n117 VDD.n116 57.1093
R4826 VDD.n299 VDD.n52 57.1093
R4827 VDD.n135 VDD.n117 56.1076
R4828 VDD.n141 VDD.n117 56.1076
R4829 VDD.n133 VDD.n117 56.1076
R4830 VDD.n148 VDD.n117 56.1076
R4831 VDD.n130 VDD.n117 56.1076
R4832 VDD.n155 VDD.n117 56.1076
R4833 VDD.n162 VDD.n117 56.1076
R4834 VDD.n124 VDD.n117 56.1076
R4835 VDD.n121 VDD.n117 56.1076
R4836 VDD.n176 VDD.n117 56.1076
R4837 VDD.n179 VDD.n117 56.1076
R4838 VDD.n299 VDD.n298 56.1076
R4839 VDD.n299 VDD.n53 56.1076
R4840 VDD.n299 VDD.n56 56.1076
R4841 VDD.n300 VDD.n299 56.1076
R4842 VDD.n299 VDD.n57 56.1076
R4843 VDD.n299 VDD.n58 56.1076
R4844 VDD.n299 VDD.n59 56.1076
R4845 VDD.n299 VDD.n60 56.1076
R4846 VDD.n299 VDD.n61 56.1076
R4847 VDD.n299 VDD.n63 56.1076
R4848 VDD.n299 VDD.n64 56.1076
R4849 VDD.n159 VDD.n158 54.9652
R4850 VDD.n258 VDD.n255 54.9652
R4851 VDD.n169 VDD.n117 53.0388
R4852 VDD.n299 VDD.n62 53.0388
R4853 VDD.n0 VDD.t64 41.0864
R4854 VDD.n127 VDD.n117 38.6605
R4855 VDD.n185 VDD.n113 30.8211
R4856 VDD.n192 VDD.n191 30.8211
R4857 VDD.n198 VDD.n106 30.8211
R4858 VDD.n205 VDD.n204 30.8211
R4859 VDD.n211 VDD.n99 30.8211
R4860 VDD.n217 VDD.n92 30.8211
R4861 VDD.n223 VDD.n92 30.8211
R4862 VDD.n229 VDD.n88 30.8211
R4863 VDD.n235 VDD.n84 30.8211
R4864 VDD.n241 VDD.n80 30.8211
R4865 VDD.n247 VDD.n76 30.8211
R4866 VDD.n285 VDD.n71 30.8211
R4867 VDD.n99 VDD.t2 30.3679
R4868 VDD.t55 VDD.n88 30.3679
R4869 VDD.n204 VDD.t0 29.4614
R4870 VDD.t4 VDD.n84 29.4614
R4871 VDD.n167 VDD.n120 29.3652
R4872 VDD.n146 VDD.n145 29.3652
R4873 VDD.n54 VDD.n48 29.3652
R4874 VDD.n271 VDD.n270 29.3652
R4875 VDD.n8 VDD.t61 28.5655
R4876 VDD.n8 VDD.t70 28.5655
R4877 VDD.n6 VDD.t57 28.5655
R4878 VDD.n6 VDD.t53 28.5655
R4879 VDD.n4 VDD.t66 28.5655
R4880 VDD.n4 VDD.t63 28.5655
R4881 VDD.n2 VDD.t59 28.5655
R4882 VDD.n2 VDD.t69 28.5655
R4883 VDD.t29 VDD.n42 28.5655
R4884 VDD.n42 VDD.t32 28.5655
R4885 VDD.t32 VDD.n41 28.5655
R4886 VDD.n41 VDD.t8 28.5655
R4887 VDD.t50 VDD.n43 28.5655
R4888 VDD.n43 VDD.t29 28.5655
R4889 VDD.n44 VDD.t5 28.5655
R4890 VDD.n44 VDD.t50 28.5655
R4891 VDD.n27 VDD.t3 28.5655
R4892 VDD.n27 VDD.t76 28.5655
R4893 VDD.n23 VDD.t12 28.5655
R4894 VDD.t48 VDD.n23 28.5655
R4895 VDD.n14 VDD.t36 28.5655
R4896 VDD.n14 VDD.t12 28.5655
R4897 VDD.n24 VDD.t48 28.5655
R4898 VDD.t26 VDD.n24 28.5655
R4899 VDD.n25 VDD.t26 28.5655
R4900 VDD.n25 VDD.t1 28.5655
R4901 VDD.n340 VDD.t73 28.5655
R4902 VDD.n340 VDD.t15 28.5655
R4903 VDD.t38 VDD.n338 28.5655
R4904 VDD.n338 VDD.t43 28.5655
R4905 VDD.t43 VDD.n337 28.5655
R4906 VDD.n337 VDD.t20 28.5655
R4907 VDD.t15 VDD.n339 28.5655
R4908 VDD.n339 VDD.t38 28.5655
R4909 VDD.n321 VDD.t34 28.5655
R4910 VDD.n321 VDD.t74 28.5655
R4911 VDD.n319 VDD.t23 28.5655
R4912 VDD.t52 VDD.n319 28.5655
R4913 VDD.n310 VDD.t45 28.5655
R4914 VDD.n310 VDD.t23 28.5655
R4915 VDD.n320 VDD.t52 28.5655
R4916 VDD.t34 VDD.n320 28.5655
R4917 VDD.n323 VDD.t75 28.5655
R4918 VDD.n323 VDD.t72 28.5655
R4919 VDD.n350 VDD.t54 28.5655
R4920 VDD.n350 VDD.t40 28.5655
R4921 VDD.n348 VDD.t60 28.5655
R4922 VDD.n348 VDD.t68 28.5655
R4923 VDD.n346 VDD.t56 28.5655
R4924 VDD.n346 VDD.t71 28.5655
R4925 VDD.n344 VDD.t65 28.5655
R4926 VDD.n344 VDD.t62 28.5655
R4927 VDD.n343 VDD.t58 28.5655
R4928 VDD.n343 VDD.t67 28.5655
R4929 VDD.n106 VDD.t25 28.5549
R4930 VDD.t14 VDD.n80 28.5549
R4931 VDD.n191 VDD.t47 27.6484
R4932 VDD.t28 VDD.n76 27.6484
R4933 VDD.n113 VDD.t11 26.7419
R4934 VDD.t31 VDD.n71 26.7419
R4935 VDD.n116 VDD.t17 25.8354
R4936 VDD.t7 VDD.n52 25.8354
R4937 VDD.n183 VDD.n182 25.6005
R4938 VDD.n183 VDD.n108 25.6005
R4939 VDD.n194 VDD.n108 25.6005
R4940 VDD.n195 VDD.n194 25.6005
R4941 VDD.n196 VDD.n195 25.6005
R4942 VDD.n196 VDD.n101 25.6005
R4943 VDD.n207 VDD.n101 25.6005
R4944 VDD.n208 VDD.n207 25.6005
R4945 VDD.n209 VDD.n208 25.6005
R4946 VDD.n209 VDD.n94 25.6005
R4947 VDD.n219 VDD.n94 25.6005
R4948 VDD.n220 VDD.n219 25.6005
R4949 VDD.n221 VDD.n220 25.6005
R4950 VDD.n221 VDD.n86 25.6005
R4951 VDD.n231 VDD.n86 25.6005
R4952 VDD.n232 VDD.n231 25.6005
R4953 VDD.n233 VDD.n232 25.6005
R4954 VDD.n233 VDD.n78 25.6005
R4955 VDD.n243 VDD.n78 25.6005
R4956 VDD.n244 VDD.n243 25.6005
R4957 VDD.n245 VDD.n244 25.6005
R4958 VDD.n245 VDD.n69 25.6005
R4959 VDD.n287 VDD.n69 25.6005
R4960 VDD.n288 VDD.n287 25.6005
R4961 VDD.n181 VDD.n115 25.6005
R4962 VDD.n118 VDD.n115 25.6005
R4963 VDD.n174 VDD.n118 25.6005
R4964 VDD.n174 VDD.n173 25.6005
R4965 VDD.n173 VDD.n172 25.6005
R4966 VDD.n172 VDD.n120 25.6005
R4967 VDD.n167 VDD.n166 25.6005
R4968 VDD.n166 VDD.n165 25.6005
R4969 VDD.n165 VDD.n123 25.6005
R4970 VDD.n160 VDD.n123 25.6005
R4971 VDD.n160 VDD.n159 25.6005
R4972 VDD.n158 VDD.n126 25.6005
R4973 VDD.n153 VDD.n126 25.6005
R4974 VDD.n153 VDD.n152 25.6005
R4975 VDD.n152 VDD.n151 25.6005
R4976 VDD.n151 VDD.n129 25.6005
R4977 VDD.n146 VDD.n129 25.6005
R4978 VDD.n145 VDD.n144 25.6005
R4979 VDD.n144 VDD.n132 25.6005
R4980 VDD.n139 VDD.n132 25.6005
R4981 VDD.n139 VDD.n138 25.6005
R4982 VDD.n138 VDD.n137 25.6005
R4983 VDD.n187 VDD.n111 25.6005
R4984 VDD.n188 VDD.n187 25.6005
R4985 VDD.n189 VDD.n188 25.6005
R4986 VDD.n189 VDD.n104 25.6005
R4987 VDD.n200 VDD.n104 25.6005
R4988 VDD.n201 VDD.n200 25.6005
R4989 VDD.n202 VDD.n201 25.6005
R4990 VDD.n202 VDD.n97 25.6005
R4991 VDD.n213 VDD.n97 25.6005
R4992 VDD.n214 VDD.n213 25.6005
R4993 VDD.n215 VDD.n214 25.6005
R4994 VDD.n215 VDD.n90 25.6005
R4995 VDD.n225 VDD.n90 25.6005
R4996 VDD.n226 VDD.n225 25.6005
R4997 VDD.n227 VDD.n226 25.6005
R4998 VDD.n227 VDD.n82 25.6005
R4999 VDD.n237 VDD.n82 25.6005
R5000 VDD.n238 VDD.n237 25.6005
R5001 VDD.n239 VDD.n238 25.6005
R5002 VDD.n239 VDD.n74 25.6005
R5003 VDD.n249 VDD.n74 25.6005
R5004 VDD.n250 VDD.n249 25.6005
R5005 VDD.n283 VDD.n250 25.6005
R5006 VDD.n283 VDD.n282 25.6005
R5007 VDD.n296 VDD.n295 25.6005
R5008 VDD.n295 VDD.n294 25.6005
R5009 VDD.n294 VDD.n293 25.6005
R5010 VDD.n293 VDD.n291 25.6005
R5011 VDD.n291 VDD.n47 25.6005
R5012 VDD.n54 VDD.n47 25.6005
R5013 VDD.n302 VDD.n49 25.6005
R5014 VDD.n251 VDD.n49 25.6005
R5015 VDD.n254 VDD.n251 25.6005
R5016 VDD.n255 VDD.n254 25.6005
R5017 VDD.n259 VDD.n258 25.6005
R5018 VDD.n262 VDD.n259 25.6005
R5019 VDD.n263 VDD.n262 25.6005
R5020 VDD.n266 VDD.n263 25.6005
R5021 VDD.n267 VDD.n266 25.6005
R5022 VDD.n270 VDD.n267 25.6005
R5023 VDD.n274 VDD.n271 25.6005
R5024 VDD.n275 VDD.n274 25.6005
R5025 VDD.n278 VDD.n275 25.6005
R5026 VDD.n280 VDD.n278 25.6005
R5027 VDD.n281 VDD.n280 25.6005
R5028 VDD.n303 VDD.n302 23.3417
R5029 VDD.n0 VDD.t18 14.285
R5030 VDD.n304 VDD.n303 9.3686
R5031 VDD.n304 VDD.n47 9.36343
R5032 VDD.n185 VDD.t17 4.98619
R5033 VDD.n285 VDD.t7 4.98619
R5034 VDD.n192 VDD.t11 4.0797
R5035 VDD.n247 VDD.t31 4.0797
R5036 VDD.n28 VDD.n26 3.35217
R5037 VDD.n324 VDD.n322 3.35217
R5038 VDD.n198 VDD.t47 3.17321
R5039 VDD.n241 VDD.t28 3.17321
R5040 VDD.n3 VDD.n1 3.06997
R5041 VDD.n46 VDD.n45 2.73818
R5042 VDD.n342 VDD.n341 2.73818
R5043 VDD VDD.n356 2.6239
R5044 VDD.n353 VDD.n352 2.45598
R5045 VDD.n205 VDD.t25 2.26672
R5046 VDD.n235 VDD.t14 2.26672
R5047 VDD.n303 VDD.n48 2.25932
R5048 VDD.n305 VDD.n304 2.20937
R5049 VDD.n354 VDD.n342 2.07758
R5050 VDD.n356 VDD.n9 1.76955
R5051 VDD.n354 VDD.n353 1.63948
R5052 VDD.n305 VDD.n46 1.485
R5053 VDD.n211 VDD.t0 1.36023
R5054 VDD.n229 VDD.t4 1.36023
R5055 VDD.n355 VDD.n354 0.9725
R5056 VDD.n5 VDD.n3 0.61449
R5057 VDD.n7 VDD.n5 0.61449
R5058 VDD.n9 VDD.n7 0.61449
R5059 VDD.n46 VDD.n28 0.61449
R5060 VDD.n342 VDD.n324 0.61449
R5061 VDD.n347 VDD.n345 0.61449
R5062 VDD.n349 VDD.n347 0.61449
R5063 VDD.n353 VDD.n349 0.61449
R5064 VDD.n355 VDD.n305 0.590949
R5065 VDD.n356 VDD.n355 0.4865
R5066 VDD.n217 VDD.t2 0.453744
R5067 VDD.n223 VDD.t55 0.453744
R5068 VDD.n336 VDD.n327 0.38373
R5069 VDD.n331 VDD.n326 0.38373
R5070 VDD.n312 VDD.n311 0.38373
R5071 VDD.n318 VDD.n307 0.38373
R5072 VDD.n40 VDD.n39 0.383729
R5073 VDD.n33 VDD.n30 0.383729
R5074 VDD.n15 VDD.n13 0.383729
R5075 VDD.n22 VDD.n21 0.383729
R5076 VDD.n35 VDD.n31 0.338735
R5077 VDD.n35 VDD.n29 0.338735
R5078 VDD.n45 VDD.n29 0.338735
R5079 VDD.n16 VDD.n11 0.338735
R5080 VDD.n11 VDD.n10 0.338735
R5081 VDD.n26 VDD.n10 0.338735
R5082 VDD.n335 VDD.n328 0.338735
R5083 VDD.n328 VDD.n325 0.338735
R5084 VDD.n341 VDD.n325 0.338735
R5085 VDD.n317 VDD.n308 0.338735
R5086 VDD.n317 VDD.n306 0.338735
R5087 VDD.n322 VDD.n306 0.338735
R5088 VDD.n38 VDD.n31 0.285826
R5089 VDD.n36 VDD.n35 0.285826
R5090 VDD.n17 VDD.n16 0.285826
R5091 VDD.n19 VDD.n11 0.285826
R5092 VDD.n335 VDD.n334 0.285826
R5093 VDD.n329 VDD.n328 0.285826
R5094 VDD.n309 VDD.n308 0.285826
R5095 VDD.n317 VDD.n316 0.285826
R5096 VDD.n37 VDD.n36 0.188
R5097 VDD.n38 VDD.n37 0.188
R5098 VDD.n34 VDD.n33 0.188
R5099 VDD.n33 VDD.n32 0.188
R5100 VDD.n39 VDD.n32 0.188
R5101 VDD.n18 VDD.n17 0.188
R5102 VDD.n19 VDD.n18 0.188
R5103 VDD.n13 VDD.n12 0.188
R5104 VDD.n21 VDD.n12 0.188
R5105 VDD.n21 VDD.n20 0.188
R5106 VDD.n331 VDD.n330 0.188
R5107 VDD.n332 VDD.n331 0.188
R5108 VDD.n332 VDD.n327 0.188
R5109 VDD.n333 VDD.n329 0.188
R5110 VDD.n334 VDD.n333 0.188
R5111 VDD.n313 VDD.n312 0.188
R5112 VDD.n313 VDD.n307 0.188
R5113 VDD.n315 VDD.n307 0.188
R5114 VDD.n314 VDD.n309 0.188
R5115 VDD.n316 VDD.n314 0.188
R5116 VDD.n40 VDD.n31 0.0984044
R5117 VDD.n35 VDD.n30 0.0984044
R5118 VDD.n16 VDD.n15 0.0984044
R5119 VDD.n22 VDD.n11 0.0984044
R5120 VDD.n328 VDD.n326 0.0984028
R5121 VDD.n336 VDD.n335 0.0984028
R5122 VDD.n318 VDD.n317 0.0984028
R5123 VDD.n311 VDD.n308 0.0984028
R5124 VDD.n352 VDD.n351 0.0793043
R5125 a_2080_2896.n68 a_2080_2896.n67 185
R5126 a_2080_2896.n68 a_2080_2896.n55 185
R5127 a_2080_2896.n68 a_2080_2896.n54 185
R5128 a_2080_2896.n68 a_2080_2896.n52 185
R5129 a_2080_2896.n68 a_2080_2896.n51 185
R5130 a_2080_2896.n69 a_2080_2896.n68 185
R5131 a_2080_2896.n91 a_2080_2896.n5 185
R5132 a_2080_2896.n91 a_2080_2896.n3 185
R5133 a_2080_2896.n91 a_2080_2896.n6 185
R5134 a_2080_2896.n91 a_2080_2896.n2 185
R5135 a_2080_2896.n91 a_2080_2896.n7 185
R5136 a_2080_2896.n91 a_2080_2896.n1 185
R5137 a_2080_2896.n91 a_2080_2896.n90 185
R5138 a_2080_2896.n36 a_2080_2896.t35 165.607
R5139 a_2080_2896.n24 a_2080_2896.t22 165.607
R5140 a_2080_2896.n85 a_2080_2896.t20 165.032
R5141 a_2080_2896.n34 a_2080_2896.t21 165.032
R5142 a_2080_2896.n33 a_2080_2896.t8 165.032
R5143 a_2080_2896.n32 a_2080_2896.t18 165.032
R5144 a_2080_2896.n31 a_2080_2896.t29 165.032
R5145 a_2080_2896.n30 a_2080_2896.t28 165.032
R5146 a_2080_2896.n29 a_2080_2896.t39 165.032
R5147 a_2080_2896.n28 a_2080_2896.t40 165.032
R5148 a_2080_2896.n27 a_2080_2896.t11 165.032
R5149 a_2080_2896.n26 a_2080_2896.t10 165.032
R5150 a_2080_2896.n25 a_2080_2896.t9 165.032
R5151 a_2080_2896.n24 a_2080_2896.t30 165.032
R5152 a_2080_2896.n83 a_2080_2896.t42 163.058
R5153 a_2080_2896.n81 a_2080_2896.t31 163.058
R5154 a_2080_2896.n79 a_2080_2896.t41 163.058
R5155 a_2080_2896.n77 a_2080_2896.t13 163.058
R5156 a_2080_2896.n75 a_2080_2896.t12 163.058
R5157 a_2080_2896.n47 a_2080_2896.t25 163.058
R5158 a_2080_2896.n73 a_2080_2896.t23 163.058
R5159 a_2080_2896.n43 a_2080_2896.t34 163.058
R5160 a_2080_2896.n41 a_2080_2896.t33 163.058
R5161 a_2080_2896.n39 a_2080_2896.t32 163.058
R5162 a_2080_2896.n37 a_2080_2896.t15 163.058
R5163 a_2080_2896.n35 a_2080_2896.t43 163.058
R5164 a_2080_2896.t4 a_2080_2896.n71 162.941
R5165 a_2080_2896.n71 a_2080_2896.t6 162.941
R5166 a_2080_2896.n83 a_2080_2896.t26 162.781
R5167 a_2080_2896.n81 a_2080_2896.t14 162.781
R5168 a_2080_2896.n79 a_2080_2896.t24 162.781
R5169 a_2080_2896.n77 a_2080_2896.t37 162.781
R5170 a_2080_2896.n75 a_2080_2896.t36 162.781
R5171 a_2080_2896.n43 a_2080_2896.t19 162.781
R5172 a_2080_2896.n41 a_2080_2896.t17 162.781
R5173 a_2080_2896.n39 a_2080_2896.t16 162.781
R5174 a_2080_2896.n37 a_2080_2896.t38 162.781
R5175 a_2080_2896.n35 a_2080_2896.t27 162.781
R5176 a_2080_2896.n72 a_2080_2896.t4 162.639
R5177 a_2080_2896.t6 a_2080_2896.n48 162.639
R5178 a_2080_2896.n9 a_2080_2896.t1 130.75
R5179 a_2080_2896.n9 a_2080_2896.t3 91.3557
R5180 a_2080_2896.n68 a_2080_2896.n53 86.5152
R5181 a_2080_2896.n91 a_2080_2896.n0 86.5152
R5182 a_2080_2896.n11 a_2080_2896.n4 30.3012
R5183 a_2080_2896.n61 a_2080_2896.n54 24.8476
R5184 a_2080_2896.n59 a_2080_2896.n52 24.8476
R5185 a_2080_2896.n90 a_2080_2896.n89 24.8476
R5186 a_2080_2896.n63 a_2080_2896.n55 23.3417
R5187 a_2080_2896.n57 a_2080_2896.n51 23.3417
R5188 a_2080_2896.n8 a_2080_2896.n1 23.3417
R5189 a_2080_2896.n87 a_2080_2896.n0 22.0256
R5190 a_2080_2896.n67 a_2080_2896.n66 21.8358
R5191 a_2080_2896.n69 a_2080_2896.n50 21.8358
R5192 a_2080_2896.n21 a_2080_2896.n7 21.8358
R5193 a_2080_2896.n19 a_2080_2896.n2 20.3299
R5194 a_2080_2896.n17 a_2080_2896.n6 18.824
R5195 a_2080_2896.n15 a_2080_2896.n3 17.3181
R5196 a_2080_2896.n91 a_2080_2896.n4 16.3559
R5197 a_2080_2896.n13 a_2080_2896.n5 15.8123
R5198 a_2080_2896.n67 a_2080_2896.n56 14.5711
R5199 a_2080_2896.n70 a_2080_2896.n69 14.5711
R5200 a_2080_2896.n87 a_2080_2896.n86 12.9589
R5201 a_2080_2896.n61 a_2080_2896.n53 12.7256
R5202 a_2080_2896.n59 a_2080_2896.n53 12.7256
R5203 a_2080_2896.n89 a_2080_2896.n0 12.7256
R5204 a_2080_2896.n11 a_2080_2896.n5 11.2946
R5205 a_2080_2896.n13 a_2080_2896.n3 9.78874
R5206 a_2080_2896.n62 a_2080_2896.n61 9.3005
R5207 a_2080_2896.n64 a_2080_2896.n63 9.3005
R5208 a_2080_2896.n66 a_2080_2896.n65 9.3005
R5209 a_2080_2896.n60 a_2080_2896.n59 9.3005
R5210 a_2080_2896.n58 a_2080_2896.n57 9.3005
R5211 a_2080_2896.n50 a_2080_2896.n49 9.3005
R5212 a_2080_2896.n89 a_2080_2896.n88 9.3005
R5213 a_2080_2896.n23 a_2080_2896.n8 9.3005
R5214 a_2080_2896.n22 a_2080_2896.n21 9.3005
R5215 a_2080_2896.n20 a_2080_2896.n19 9.3005
R5216 a_2080_2896.n18 a_2080_2896.n17 9.3005
R5217 a_2080_2896.n16 a_2080_2896.n15 9.3005
R5218 a_2080_2896.n14 a_2080_2896.n13 9.3005
R5219 a_2080_2896.n12 a_2080_2896.n11 9.3005
R5220 a_2080_2896.n86 a_2080_2896.n85 8.61608
R5221 a_2080_2896.n15 a_2080_2896.n6 8.28285
R5222 a_2080_2896.n17 a_2080_2896.n2 6.77697
R5223 a_2080_2896.n68 a_2080_2896.t7 5.8005
R5224 a_2080_2896.n68 a_2080_2896.t5 5.8005
R5225 a_2080_2896.n19 a_2080_2896.n7 5.27109
R5226 a_2080_2896.n66 a_2080_2896.n55 3.76521
R5227 a_2080_2896.n51 a_2080_2896.n50 3.76521
R5228 a_2080_2896.n21 a_2080_2896.n1 3.76521
R5229 a_2080_2896.t0 a_2080_2896.n91 2.48621
R5230 a_2080_2896.n91 a_2080_2896.t2 2.48621
R5231 a_2080_2896.n10 a_2080_2896.n4 2.36936
R5232 a_2080_2896.n63 a_2080_2896.n54 2.25932
R5233 a_2080_2896.n57 a_2080_2896.n52 2.25932
R5234 a_2080_2896.n90 a_2080_2896.n8 2.25932
R5235 a_2080_2896.n84 a_2080_2896.n83 2.25162
R5236 a_2080_2896.n82 a_2080_2896.n81 2.25162
R5237 a_2080_2896.n80 a_2080_2896.n79 2.25162
R5238 a_2080_2896.n78 a_2080_2896.n77 2.25162
R5239 a_2080_2896.n76 a_2080_2896.n75 2.25162
R5240 a_2080_2896.n47 a_2080_2896.n45 2.25162
R5241 a_2080_2896.n74 a_2080_2896.n73 2.25162
R5242 a_2080_2896.n44 a_2080_2896.n43 2.25162
R5243 a_2080_2896.n42 a_2080_2896.n41 2.25162
R5244 a_2080_2896.n40 a_2080_2896.n39 2.25162
R5245 a_2080_2896.n38 a_2080_2896.n37 2.25162
R5246 a_2080_2896.n36 a_2080_2896.n35 2.25162
R5247 a_2080_2896.n86 a_2080_2896.n34 2.17137
R5248 a_2080_2896.n38 a_2080_2896.n36 0.574917
R5249 a_2080_2896.n40 a_2080_2896.n38 0.574917
R5250 a_2080_2896.n42 a_2080_2896.n40 0.574917
R5251 a_2080_2896.n44 a_2080_2896.n42 0.574917
R5252 a_2080_2896.n45 a_2080_2896.n44 0.574917
R5253 a_2080_2896.n74 a_2080_2896.n45 0.574917
R5254 a_2080_2896.n76 a_2080_2896.n74 0.574917
R5255 a_2080_2896.n78 a_2080_2896.n76 0.574917
R5256 a_2080_2896.n80 a_2080_2896.n78 0.574917
R5257 a_2080_2896.n82 a_2080_2896.n80 0.574917
R5258 a_2080_2896.n84 a_2080_2896.n82 0.574917
R5259 a_2080_2896.n85 a_2080_2896.n84 0.574917
R5260 a_2080_2896.n25 a_2080_2896.n24 0.574917
R5261 a_2080_2896.n26 a_2080_2896.n25 0.574917
R5262 a_2080_2896.n27 a_2080_2896.n26 0.574917
R5263 a_2080_2896.n28 a_2080_2896.n27 0.574917
R5264 a_2080_2896.n29 a_2080_2896.n28 0.574917
R5265 a_2080_2896.n30 a_2080_2896.n29 0.574917
R5266 a_2080_2896.n31 a_2080_2896.n30 0.574917
R5267 a_2080_2896.n32 a_2080_2896.n31 0.574917
R5268 a_2080_2896.n33 a_2080_2896.n32 0.574917
R5269 a_2080_2896.n34 a_2080_2896.n33 0.574917
R5270 a_2080_2896.n10 a_2080_2896.n9 0.320353
R5271 a_2080_2896.n48 a_2080_2896.n46 0.302413
R5272 a_2080_2896.n72 a_2080_2896.n46 0.302413
R5273 a_2080_2896.n56 a_2080_2896.n46 0.217891
R5274 a_2080_2896.n71 a_2080_2896.n70 0.217891
R5275 a_2080_2896.n65 a_2080_2896.n56 0.196152
R5276 a_2080_2896.n65 a_2080_2896.n64 0.196152
R5277 a_2080_2896.n64 a_2080_2896.n62 0.196152
R5278 a_2080_2896.n62 a_2080_2896.n60 0.196152
R5279 a_2080_2896.n60 a_2080_2896.n58 0.196152
R5280 a_2080_2896.n58 a_2080_2896.n49 0.196152
R5281 a_2080_2896.n70 a_2080_2896.n49 0.196152
R5282 a_2080_2896.n12 a_2080_2896.n10 0.196152
R5283 a_2080_2896.n14 a_2080_2896.n12 0.196152
R5284 a_2080_2896.n16 a_2080_2896.n14 0.196152
R5285 a_2080_2896.n18 a_2080_2896.n16 0.196152
R5286 a_2080_2896.n20 a_2080_2896.n18 0.196152
R5287 a_2080_2896.n22 a_2080_2896.n20 0.196152
R5288 a_2080_2896.n23 a_2080_2896.n22 0.196152
R5289 a_2080_2896.n88 a_2080_2896.n23 0.196152
R5290 a_2080_2896.n88 a_2080_2896.n87 0.196152
R5291 a_2080_2896.n48 a_2080_2896.n47 0.142018
R5292 a_2080_2896.n73 a_2080_2896.n72 0.142018
R5293 a_4920_2896.n46 a_4920_2896.n28 185
R5294 a_4920_2896.n46 a_4920_2896.n27 185
R5295 a_4920_2896.n46 a_4920_2896.n26 185
R5296 a_4920_2896.n46 a_4920_2896.n25 185
R5297 a_4920_2896.n46 a_4920_2896.n24 185
R5298 a_4920_2896.n46 a_4920_2896.n23 185
R5299 a_4920_2896.n46 a_4920_2896.n22 185
R5300 a_4920_2896.n30 a_4920_2896.t25 130.75
R5301 a_4920_2896.n30 a_4920_2896.t26 91.3557
R5302 a_4920_2896.n47 a_4920_2896.n46 86.5152
R5303 a_4920_2896.n45 a_4920_2896.n29 30.3012
R5304 a_4920_2896.n15 a_4920_2896.n14 26.8581
R5305 a_4920_2896.n5 a_4920_2896.n4 26.6299
R5306 a_4920_2896.n19 a_4920_2896.n9 25.7063
R5307 a_4920_2896.n18 a_4920_2896.n10 25.7063
R5308 a_4920_2896.n17 a_4920_2896.n11 25.7063
R5309 a_4920_2896.n16 a_4920_2896.n12 25.7063
R5310 a_4920_2896.n15 a_4920_2896.n13 25.7063
R5311 a_4920_2896.n51 a_4920_2896.n50 25.4783
R5312 a_4920_2896.n5 a_4920_2896.n3 25.4781
R5313 a_4920_2896.n6 a_4920_2896.n2 25.4781
R5314 a_4920_2896.n7 a_4920_2896.n1 25.4781
R5315 a_4920_2896.n8 a_4920_2896.n0 25.4781
R5316 a_4920_2896.n22 a_4920_2896.n21 24.8476
R5317 a_4920_2896.n31 a_4920_2896.n23 23.3417
R5318 a_4920_2896.n48 a_4920_2896.n47 22.0256
R5319 a_4920_2896.n33 a_4920_2896.n24 21.8358
R5320 a_4920_2896.n35 a_4920_2896.n25 20.3299
R5321 a_4920_2896.n37 a_4920_2896.n26 18.824
R5322 a_4920_2896.n39 a_4920_2896.n27 17.3181
R5323 a_4920_2896.n46 a_4920_2896.n45 16.3559
R5324 a_4920_2896.n41 a_4920_2896.n28 15.8123
R5325 a_4920_2896.n47 a_4920_2896.n21 12.7256
R5326 a_4920_2896.n29 a_4920_2896.n28 11.2946
R5327 a_4920_2896.n41 a_4920_2896.n27 9.78874
R5328 a_4920_2896.n49 a_4920_2896.n19 9.30285
R5329 a_4920_2896.n21 a_4920_2896.n20 9.3005
R5330 a_4920_2896.n32 a_4920_2896.n31 9.3005
R5331 a_4920_2896.n34 a_4920_2896.n33 9.3005
R5332 a_4920_2896.n36 a_4920_2896.n35 9.3005
R5333 a_4920_2896.n38 a_4920_2896.n37 9.3005
R5334 a_4920_2896.n40 a_4920_2896.n39 9.3005
R5335 a_4920_2896.n42 a_4920_2896.n41 9.3005
R5336 a_4920_2896.n43 a_4920_2896.n29 9.3005
R5337 a_4920_2896.n39 a_4920_2896.n26 8.28285
R5338 a_4920_2896.n37 a_4920_2896.n25 6.77697
R5339 a_4920_2896.n4 a_4920_2896.t14 5.8005
R5340 a_4920_2896.n4 a_4920_2896.t9 5.8005
R5341 a_4920_2896.n3 a_4920_2896.t22 5.8005
R5342 a_4920_2896.n3 a_4920_2896.t21 5.8005
R5343 a_4920_2896.n2 a_4920_2896.t20 5.8005
R5344 a_4920_2896.n2 a_4920_2896.t3 5.8005
R5345 a_4920_2896.n1 a_4920_2896.t4 5.8005
R5346 a_4920_2896.n1 a_4920_2896.t11 5.8005
R5347 a_4920_2896.n0 a_4920_2896.t10 5.8005
R5348 a_4920_2896.n0 a_4920_2896.t16 5.8005
R5349 a_4920_2896.n9 a_4920_2896.t8 5.8005
R5350 a_4920_2896.n9 a_4920_2896.t1 5.8005
R5351 a_4920_2896.n10 a_4920_2896.t18 5.8005
R5352 a_4920_2896.n10 a_4920_2896.t2 5.8005
R5353 a_4920_2896.n11 a_4920_2896.t13 5.8005
R5354 a_4920_2896.n11 a_4920_2896.t19 5.8005
R5355 a_4920_2896.n12 a_4920_2896.t5 5.8005
R5356 a_4920_2896.n12 a_4920_2896.t12 5.8005
R5357 a_4920_2896.n13 a_4920_2896.t7 5.8005
R5358 a_4920_2896.n13 a_4920_2896.t6 5.8005
R5359 a_4920_2896.n14 a_4920_2896.t0 5.8005
R5360 a_4920_2896.n14 a_4920_2896.t17 5.8005
R5361 a_4920_2896.t23 a_4920_2896.n51 5.8005
R5362 a_4920_2896.n51 a_4920_2896.t15 5.8005
R5363 a_4920_2896.n35 a_4920_2896.n24 5.27109
R5364 a_4920_2896.n33 a_4920_2896.n23 3.76521
R5365 a_4920_2896.n50 a_4920_2896.n49 2.92217
R5366 a_4920_2896.n46 a_4920_2896.t26 2.48621
R5367 a_4920_2896.n46 a_4920_2896.t24 2.48621
R5368 a_4920_2896.n45 a_4920_2896.n44 2.36936
R5369 a_4920_2896.n31 a_4920_2896.n22 2.25932
R5370 a_4920_2896.n49 a_4920_2896.n48 2.19829
R5371 a_4920_2896.n16 a_4920_2896.n15 1.15229
R5372 a_4920_2896.n17 a_4920_2896.n16 1.15229
R5373 a_4920_2896.n18 a_4920_2896.n17 1.15229
R5374 a_4920_2896.n19 a_4920_2896.n18 1.15229
R5375 a_4920_2896.n6 a_4920_2896.n5 1.15229
R5376 a_4920_2896.n7 a_4920_2896.n6 1.15229
R5377 a_4920_2896.n8 a_4920_2896.n7 1.15229
R5378 a_4920_2896.n50 a_4920_2896.n8 1.15229
R5379 a_4920_2896.n44 a_4920_2896.n30 0.320353
R5380 a_4920_2896.n44 a_4920_2896.n43 0.196152
R5381 a_4920_2896.n43 a_4920_2896.n42 0.196152
R5382 a_4920_2896.n42 a_4920_2896.n40 0.196152
R5383 a_4920_2896.n40 a_4920_2896.n38 0.196152
R5384 a_4920_2896.n38 a_4920_2896.n36 0.196152
R5385 a_4920_2896.n36 a_4920_2896.n34 0.196152
R5386 a_4920_2896.n34 a_4920_2896.n32 0.196152
R5387 a_4920_2896.n32 a_4920_2896.n20 0.196152
R5388 a_4920_2896.n48 a_4920_2896.n20 0.196152
R5389 VP.n0 VP.t7 263.647
R5390 VP.n3 VP.t3 262.863
R5391 VP.n2 VP.t1 262.498
R5392 VP.n0 VP.t6 261.709
R5393 VP.n1 VP.t2 261.709
R5394 VP.n3 VP.t5 261.584
R5395 VP.n4 VP.t4 261.584
R5396 VP.n5 VP.t0 261.433
R5397 VP.n6 VP.n2 8.91142
R5398 VP VP.n6 2.39915
R5399 VP.n1 VP.n0 1.72698
R5400 VP.n6 VP.n5 1.52193
R5401 VP.n5 VP.n4 1.4312
R5402 VP.n4 VP.n3 1.16675
R5403 VP.n2 VP.n1 1.14999
R5404 a_2995_7336.n30 a_2995_7336.n29 185
R5405 a_2995_7336.n30 a_2995_7336.n12 185
R5406 a_2995_7336.n30 a_2995_7336.n11 185
R5407 a_2995_7336.n30 a_2995_7336.n10 185
R5408 a_2995_7336.n30 a_2995_7336.n9 185
R5409 a_2995_7336.n30 a_2995_7336.n8 185
R5410 a_2995_7336.n30 a_2995_7336.n7 185
R5411 a_2995_7336.n13 a_2995_7336.t17 130.75
R5412 a_2995_7336.n13 a_2995_7336.t19 91.3557
R5413 a_2995_7336.n31 a_2995_7336.n30 86.5152
R5414 a_2995_7336.n15 a_2995_7336.n6 30.3012
R5415 a_2995_7336.n29 a_2995_7336.n5 24.8476
R5416 a_2995_7336.n28 a_2995_7336.n12 23.3417
R5417 a_2995_7336.n32 a_2995_7336.n31 22.0256
R5418 a_2995_7336.n25 a_2995_7336.n11 21.8358
R5419 a_2995_7336.n23 a_2995_7336.n10 20.3299
R5420 a_2995_7336.n21 a_2995_7336.n9 18.824
R5421 a_2995_7336.n19 a_2995_7336.n8 17.3181
R5422 a_2995_7336.n30 a_2995_7336.n6 16.3559
R5423 a_2995_7336.n17 a_2995_7336.n7 15.8123
R5424 a_2995_7336.n31 a_2995_7336.n5 12.7256
R5425 a_2995_7336.n39 a_2995_7336.n38 12.1709
R5426 a_2995_7336.n40 a_2995_7336.n39 12.1709
R5427 a_2995_7336.n38 a_2995_7336.n33 11.493
R5428 a_2995_7336.n37 a_2995_7336.n35 11.493
R5429 a_2995_7336.n3 a_2995_7336.n1 11.493
R5430 a_2995_7336.n40 a_2995_7336.n0 11.4929
R5431 a_2995_7336.n38 a_2995_7336.n34 11.4929
R5432 a_2995_7336.n37 a_2995_7336.n36 11.4929
R5433 a_2995_7336.n3 a_2995_7336.n2 11.4929
R5434 a_2995_7336.n41 a_2995_7336.n40 11.4929
R5435 a_2995_7336.n15 a_2995_7336.n7 11.2946
R5436 a_2995_7336.n17 a_2995_7336.n8 9.78874
R5437 a_2995_7336.n5 a_2995_7336.n4 9.3005
R5438 a_2995_7336.n28 a_2995_7336.n27 9.3005
R5439 a_2995_7336.n26 a_2995_7336.n25 9.3005
R5440 a_2995_7336.n24 a_2995_7336.n23 9.3005
R5441 a_2995_7336.n22 a_2995_7336.n21 9.3005
R5442 a_2995_7336.n20 a_2995_7336.n19 9.3005
R5443 a_2995_7336.n18 a_2995_7336.n17 9.3005
R5444 a_2995_7336.n16 a_2995_7336.n15 9.3005
R5445 a_2995_7336.n19 a_2995_7336.n9 8.28285
R5446 a_2995_7336.n21 a_2995_7336.n10 6.77697
R5447 a_2995_7336.n23 a_2995_7336.n11 5.27109
R5448 a_2995_7336.n25 a_2995_7336.n12 3.76521
R5449 a_2995_7336.n39 a_2995_7336.n32 3.48602
R5450 a_2995_7336.n0 a_2995_7336.t11 2.48621
R5451 a_2995_7336.n0 a_2995_7336.t5 2.48621
R5452 a_2995_7336.n34 a_2995_7336.t8 2.48621
R5453 a_2995_7336.n34 a_2995_7336.t13 2.48621
R5454 a_2995_7336.n33 a_2995_7336.t16 2.48621
R5455 a_2995_7336.n33 a_2995_7336.t7 2.48621
R5456 a_2995_7336.n36 a_2995_7336.t10 2.48621
R5457 a_2995_7336.n36 a_2995_7336.t4 2.48621
R5458 a_2995_7336.n35 a_2995_7336.t6 2.48621
R5459 a_2995_7336.n35 a_2995_7336.t12 2.48621
R5460 a_2995_7336.n2 a_2995_7336.t3 2.48621
R5461 a_2995_7336.n2 a_2995_7336.t15 2.48621
R5462 a_2995_7336.n1 a_2995_7336.t9 2.48621
R5463 a_2995_7336.n1 a_2995_7336.t2 2.48621
R5464 a_2995_7336.n30 a_2995_7336.t14 2.48621
R5465 a_2995_7336.n30 a_2995_7336.t18 2.48621
R5466 a_2995_7336.n41 a_2995_7336.t1 2.48621
R5467 a_2995_7336.t0 a_2995_7336.n41 2.48621
R5468 a_2995_7336.n14 a_2995_7336.n6 2.36936
R5469 a_2995_7336.n29 a_2995_7336.n28 2.25932
R5470 a_2995_7336.n38 a_2995_7336.n37 1.15229
R5471 a_2995_7336.n37 a_2995_7336.n3 1.15229
R5472 a_2995_7336.n40 a_2995_7336.n3 1.15229
R5473 a_2995_7336.n14 a_2995_7336.n13 0.320353
R5474 a_2995_7336.n32 a_2995_7336.n4 0.196152
R5475 a_2995_7336.n27 a_2995_7336.n4 0.196152
R5476 a_2995_7336.n27 a_2995_7336.n26 0.196152
R5477 a_2995_7336.n26 a_2995_7336.n24 0.196152
R5478 a_2995_7336.n24 a_2995_7336.n22 0.196152
R5479 a_2995_7336.n22 a_2995_7336.n20 0.196152
R5480 a_2995_7336.n20 a_2995_7336.n18 0.196152
R5481 a_2995_7336.n18 a_2995_7336.n16 0.196152
R5482 a_2995_7336.n16 a_2995_7336.n14 0.196152
R5483 VN.n0 VN.t0 263.647
R5484 VN.n3 VN.t2 262.863
R5485 VN.n2 VN.t5 262.498
R5486 VN.n1 VN.t4 261.709
R5487 VN.n0 VN.t1 261.709
R5488 VN.n4 VN.t7 261.584
R5489 VN.n3 VN.t6 261.584
R5490 VN.n5 VN.t3 261.433
R5491 VN.n6 VN.n2 8.91142
R5492 VN VN.n6 2.48969
R5493 VN.n1 VN.n0 1.72698
R5494 VN.n6 VN.n5 1.52193
R5495 VN.n5 VN.n4 1.4312
R5496 VN.n4 VN.n3 1.16675
R5497 VN.n2 VN.n1 1.14999
R5498 a_2479_9004.n17 a_2479_9004.t22 260.111
R5499 a_2479_9004.n15 a_2479_9004.t21 260.111
R5500 a_2479_9004.n14 a_2479_9004.t5 260.111
R5501 a_2479_9004.n12 a_2479_9004.t7 260.111
R5502 a_2479_9004.n17 a_2479_9004.t9 260.111
R5503 a_2479_9004.n15 a_2479_9004.t11 260.111
R5504 a_2479_9004.n14 a_2479_9004.t24 260.111
R5505 a_2479_9004.n12 a_2479_9004.t23 260.111
R5506 a_2479_9004.n13 a_2479_9004.n11 203.413
R5507 a_2479_9004.n16 a_2479_9004.n10 203.413
R5508 a_2479_9004.n48 a_2479_9004.n47 185
R5509 a_2479_9004.n48 a_2479_9004.n30 185
R5510 a_2479_9004.n48 a_2479_9004.n29 185
R5511 a_2479_9004.n48 a_2479_9004.n28 185
R5512 a_2479_9004.n48 a_2479_9004.n27 185
R5513 a_2479_9004.n48 a_2479_9004.n26 185
R5514 a_2479_9004.n48 a_2479_9004.n25 185
R5515 a_2479_9004.n72 a_2479_9004.n4 185
R5516 a_2479_9004.n72 a_2479_9004.n6 185
R5517 a_2479_9004.n72 a_2479_9004.n3 185
R5518 a_2479_9004.n72 a_2479_9004.n7 185
R5519 a_2479_9004.n72 a_2479_9004.n2 185
R5520 a_2479_9004.n72 a_2479_9004.n8 185
R5521 a_2479_9004.n72 a_2479_9004.n1 185
R5522 a_2479_9004.n0 a_2479_9004.t3 130.75
R5523 a_2479_9004.n31 a_2479_9004.t0 130.75
R5524 a_2479_9004.t4 a_2479_9004.n0 91.3557
R5525 a_2479_9004.n31 a_2479_9004.t2 91.3557
R5526 a_2479_9004.n49 a_2479_9004.n48 86.5152
R5527 a_2479_9004.n72 a_2479_9004.n5 86.5152
R5528 a_2479_9004.n33 a_2479_9004.n24 30.3012
R5529 a_2479_9004.n71 a_2479_9004.n70 30.3012
R5530 a_2479_9004.n11 a_2479_9004.t8 28.5655
R5531 a_2479_9004.n11 a_2479_9004.t6 28.5655
R5532 a_2479_9004.n10 a_2479_9004.t12 28.5655
R5533 a_2479_9004.n10 a_2479_9004.t10 28.5655
R5534 a_2479_9004.n47 a_2479_9004.n23 24.8476
R5535 a_2479_9004.n55 a_2479_9004.n4 24.8476
R5536 a_2479_9004.n46 a_2479_9004.n30 23.3417
R5537 a_2479_9004.n57 a_2479_9004.n6 23.3417
R5538 a_2479_9004.n50 a_2479_9004.n49 22.0256
R5539 a_2479_9004.n54 a_2479_9004.n5 22.0256
R5540 a_2479_9004.n43 a_2479_9004.n29 21.8358
R5541 a_2479_9004.n59 a_2479_9004.n3 21.8358
R5542 a_2479_9004.n41 a_2479_9004.n28 20.3299
R5543 a_2479_9004.n61 a_2479_9004.n7 20.3299
R5544 a_2479_9004.n39 a_2479_9004.n27 18.824
R5545 a_2479_9004.n63 a_2479_9004.n2 18.824
R5546 a_2479_9004.n20 a_2479_9004.n18 17.4823
R5547 a_2479_9004.n37 a_2479_9004.n26 17.3181
R5548 a_2479_9004.n65 a_2479_9004.n8 17.3181
R5549 a_2479_9004.n48 a_2479_9004.n24 16.3559
R5550 a_2479_9004.n72 a_2479_9004.n71 16.3559
R5551 a_2479_9004.n35 a_2479_9004.n25 15.8123
R5552 a_2479_9004.n67 a_2479_9004.n1 15.8123
R5553 a_2479_9004.n20 a_2479_9004.n19 14.6053
R5554 a_2479_9004.n52 a_2479_9004.n51 14.377
R5555 a_2479_9004.n49 a_2479_9004.n23 12.7256
R5556 a_2479_9004.n55 a_2479_9004.n5 12.7256
R5557 a_2479_9004.n33 a_2479_9004.n25 11.2946
R5558 a_2479_9004.n70 a_2479_9004.n1 11.2946
R5559 a_2479_9004.n21 a_2479_9004.n20 10.4849
R5560 a_2479_9004.n35 a_2479_9004.n26 9.78874
R5561 a_2479_9004.n67 a_2479_9004.n8 9.78874
R5562 a_2479_9004.n23 a_2479_9004.n22 9.3005
R5563 a_2479_9004.n46 a_2479_9004.n45 9.3005
R5564 a_2479_9004.n44 a_2479_9004.n43 9.3005
R5565 a_2479_9004.n42 a_2479_9004.n41 9.3005
R5566 a_2479_9004.n40 a_2479_9004.n39 9.3005
R5567 a_2479_9004.n38 a_2479_9004.n37 9.3005
R5568 a_2479_9004.n36 a_2479_9004.n35 9.3005
R5569 a_2479_9004.n34 a_2479_9004.n33 9.3005
R5570 a_2479_9004.n56 a_2479_9004.n55 9.3005
R5571 a_2479_9004.n58 a_2479_9004.n57 9.3005
R5572 a_2479_9004.n60 a_2479_9004.n59 9.3005
R5573 a_2479_9004.n62 a_2479_9004.n61 9.3005
R5574 a_2479_9004.n64 a_2479_9004.n63 9.3005
R5575 a_2479_9004.n66 a_2479_9004.n65 9.3005
R5576 a_2479_9004.n68 a_2479_9004.n67 9.3005
R5577 a_2479_9004.n70 a_2479_9004.n69 9.3005
R5578 a_2479_9004.n21 a_2479_9004.n17 8.69704
R5579 a_2479_9004.n37 a_2479_9004.n27 8.28285
R5580 a_2479_9004.n65 a_2479_9004.n2 8.28285
R5581 a_2479_9004.n39 a_2479_9004.n28 6.77697
R5582 a_2479_9004.n63 a_2479_9004.n7 6.77697
R5583 a_2479_9004.n52 a_2479_9004.n50 6.19091
R5584 a_2479_9004.n41 a_2479_9004.n29 5.27109
R5585 a_2479_9004.n61 a_2479_9004.n3 5.27109
R5586 a_2479_9004.n43 a_2479_9004.n30 3.76521
R5587 a_2479_9004.n59 a_2479_9004.n6 3.76521
R5588 a_2479_9004.n54 a_2479_9004.n53 3.31388
R5589 a_2479_9004.n48 a_2479_9004.t17 2.48621
R5590 a_2479_9004.n48 a_2479_9004.t1 2.48621
R5591 a_2479_9004.n51 a_2479_9004.t14 2.48621
R5592 a_2479_9004.n51 a_2479_9004.t13 2.48621
R5593 a_2479_9004.n18 a_2479_9004.t16 2.48621
R5594 a_2479_9004.n18 a_2479_9004.t15 2.48621
R5595 a_2479_9004.n19 a_2479_9004.t20 2.48621
R5596 a_2479_9004.n19 a_2479_9004.t19 2.48621
R5597 a_2479_9004.t4 a_2479_9004.n72 2.48621
R5598 a_2479_9004.n72 a_2479_9004.t18 2.48621
R5599 a_2479_9004.n32 a_2479_9004.n24 2.36936
R5600 a_2479_9004.n71 a_2479_9004.n9 2.36936
R5601 a_2479_9004.n53 a_2479_9004.n52 2.30287
R5602 a_2479_9004.n47 a_2479_9004.n46 2.25932
R5603 a_2479_9004.n57 a_2479_9004.n4 2.25932
R5604 a_2479_9004.n53 a_2479_9004.n21 1.07418
R5605 a_2479_9004.n9 a_2479_9004.n0 0.320353
R5606 a_2479_9004.n32 a_2479_9004.n31 0.320353
R5607 a_2479_9004.n50 a_2479_9004.n22 0.196152
R5608 a_2479_9004.n45 a_2479_9004.n22 0.196152
R5609 a_2479_9004.n45 a_2479_9004.n44 0.196152
R5610 a_2479_9004.n44 a_2479_9004.n42 0.196152
R5611 a_2479_9004.n42 a_2479_9004.n40 0.196152
R5612 a_2479_9004.n40 a_2479_9004.n38 0.196152
R5613 a_2479_9004.n38 a_2479_9004.n36 0.196152
R5614 a_2479_9004.n36 a_2479_9004.n34 0.196152
R5615 a_2479_9004.n34 a_2479_9004.n32 0.196152
R5616 a_2479_9004.n56 a_2479_9004.n54 0.196152
R5617 a_2479_9004.n58 a_2479_9004.n56 0.196152
R5618 a_2479_9004.n60 a_2479_9004.n58 0.196152
R5619 a_2479_9004.n62 a_2479_9004.n60 0.196152
R5620 a_2479_9004.n64 a_2479_9004.n62 0.196152
R5621 a_2479_9004.n66 a_2479_9004.n64 0.196152
R5622 a_2479_9004.n68 a_2479_9004.n66 0.196152
R5623 a_2479_9004.n69 a_2479_9004.n68 0.196152
R5624 a_2479_9004.n69 a_2479_9004.n9 0.196152
R5625 a_2479_9004.n15 a_2479_9004.n14 0.0850588
R5626 a_2479_9004.n13 a_2479_9004.n12 0.0427794
R5627 a_2479_9004.n14 a_2479_9004.n13 0.0427794
R5628 a_2479_9004.n16 a_2479_9004.n15 0.0427794
R5629 a_2479_9004.n17 a_2479_9004.n16 0.0427794
R5630 a_3758_2896.n33 a_3758_2896.n32 185
R5631 a_3758_2896.n33 a_3758_2896.n15 185
R5632 a_3758_2896.n33 a_3758_2896.n14 185
R5633 a_3758_2896.n33 a_3758_2896.n13 185
R5634 a_3758_2896.n33 a_3758_2896.n12 185
R5635 a_3758_2896.n33 a_3758_2896.n11 185
R5636 a_3758_2896.n33 a_3758_2896.n10 185
R5637 a_3758_2896.n16 a_3758_2896.t12 130.75
R5638 a_3758_2896.n16 a_3758_2896.t13 91.3557
R5639 a_3758_2896.n34 a_3758_2896.n33 86.5152
R5640 a_3758_2896.n18 a_3758_2896.n9 30.3012
R5641 a_3758_2896.n2 a_3758_2896.n0 29.1073
R5642 a_3758_2896.n39 a_3758_2896.n38 27.9576
R5643 a_3758_2896.n37 a_3758_2896.n36 27.9576
R5644 a_3758_2896.n6 a_3758_2896.n5 27.9576
R5645 a_3758_2896.n4 a_3758_2896.n3 27.9576
R5646 a_3758_2896.n2 a_3758_2896.n1 27.9576
R5647 a_3758_2896.n32 a_3758_2896.n8 24.8476
R5648 a_3758_2896.n31 a_3758_2896.n15 23.3417
R5649 a_3758_2896.n35 a_3758_2896.n34 22.0256
R5650 a_3758_2896.n28 a_3758_2896.n14 21.8358
R5651 a_3758_2896.n26 a_3758_2896.n13 20.3299
R5652 a_3758_2896.n24 a_3758_2896.n12 18.824
R5653 a_3758_2896.n22 a_3758_2896.n11 17.3181
R5654 a_3758_2896.n33 a_3758_2896.n9 16.3559
R5655 a_3758_2896.n20 a_3758_2896.n10 15.8123
R5656 a_3758_2896.n34 a_3758_2896.n8 12.7256
R5657 a_3758_2896.n37 a_3758_2896.n35 12.0517
R5658 a_3758_2896.n18 a_3758_2896.n10 11.2946
R5659 a_3758_2896.n20 a_3758_2896.n11 9.78874
R5660 a_3758_2896.n8 a_3758_2896.n7 9.3005
R5661 a_3758_2896.n31 a_3758_2896.n30 9.3005
R5662 a_3758_2896.n29 a_3758_2896.n28 9.3005
R5663 a_3758_2896.n27 a_3758_2896.n26 9.3005
R5664 a_3758_2896.n25 a_3758_2896.n24 9.3005
R5665 a_3758_2896.n23 a_3758_2896.n22 9.3005
R5666 a_3758_2896.n21 a_3758_2896.n20 9.3005
R5667 a_3758_2896.n19 a_3758_2896.n18 9.3005
R5668 a_3758_2896.n22 a_3758_2896.n12 8.28285
R5669 a_3758_2896.n24 a_3758_2896.n13 6.77697
R5670 a_3758_2896.n36 a_3758_2896.t5 5.8005
R5671 a_3758_2896.n36 a_3758_2896.t7 5.8005
R5672 a_3758_2896.n5 a_3758_2896.t2 5.8005
R5673 a_3758_2896.n5 a_3758_2896.t1 5.8005
R5674 a_3758_2896.n3 a_3758_2896.t9 5.8005
R5675 a_3758_2896.n3 a_3758_2896.t8 5.8005
R5676 a_3758_2896.n1 a_3758_2896.t0 5.8005
R5677 a_3758_2896.n1 a_3758_2896.t10 5.8005
R5678 a_3758_2896.n0 a_3758_2896.t3 5.8005
R5679 a_3758_2896.n0 a_3758_2896.t4 5.8005
R5680 a_3758_2896.n39 a_3758_2896.t6 5.8005
R5681 a_3758_2896.t11 a_3758_2896.n39 5.8005
R5682 a_3758_2896.n26 a_3758_2896.n14 5.27109
R5683 a_3758_2896.n28 a_3758_2896.n15 3.76521
R5684 a_3758_2896.n33 a_3758_2896.t13 2.48621
R5685 a_3758_2896.n33 a_3758_2896.t14 2.48621
R5686 a_3758_2896.n17 a_3758_2896.n9 2.36936
R5687 a_3758_2896.n6 a_3758_2896.n4 2.30199
R5688 a_3758_2896.n32 a_3758_2896.n31 2.25932
R5689 a_3758_2896.n4 a_3758_2896.n2 1.1502
R5690 a_3758_2896.n38 a_3758_2896.n6 1.1502
R5691 a_3758_2896.n38 a_3758_2896.n37 1.1502
R5692 a_3758_2896.n17 a_3758_2896.n16 0.320353
R5693 a_3758_2896.n35 a_3758_2896.n7 0.196152
R5694 a_3758_2896.n30 a_3758_2896.n7 0.196152
R5695 a_3758_2896.n30 a_3758_2896.n29 0.196152
R5696 a_3758_2896.n29 a_3758_2896.n27 0.196152
R5697 a_3758_2896.n27 a_3758_2896.n25 0.196152
R5698 a_3758_2896.n25 a_3758_2896.n23 0.196152
R5699 a_3758_2896.n23 a_3758_2896.n21 0.196152
R5700 a_3758_2896.n21 a_3758_2896.n19 0.196152
R5701 a_3758_2896.n19 a_3758_2896.n17 0.196152
R5702 EN.n0 EN.t0 262.997
R5703 EN.n1 EN.t1 262.007
R5704 EN.n0 EN.t2 262.007
R5705 EN.n1 EN.n0 0.989232
R5706 EN EN.n1 0.365614
R5707 mim_cap_0.C1 mim_cap_0.C1.t0 17.4619
R5708 mim_cap_0.C1 mim_cap_0.C1.t1 0.00167066
R5709 IBIAS.n26 IBIAS.n25 185
R5710 IBIAS.n26 IBIAS.n8 185
R5711 IBIAS.n26 IBIAS.n7 185
R5712 IBIAS.n26 IBIAS.n6 185
R5713 IBIAS.n26 IBIAS.n5 185
R5714 IBIAS.n26 IBIAS.n4 185
R5715 IBIAS.n26 IBIAS.n3 185
R5716 IBIAS.n9 IBIAS.t1 130.75
R5717 IBIAS.n9 IBIAS.t2 91.3557
R5718 IBIAS.n27 IBIAS.n26 86.5152
R5719 IBIAS.n11 IBIAS.n2 30.3012
R5720 IBIAS.n25 IBIAS.n1 24.8476
R5721 IBIAS.n24 IBIAS.n8 23.3417
R5722 IBIAS.n28 IBIAS.n27 22.0256
R5723 IBIAS.n21 IBIAS.n7 21.8358
R5724 IBIAS.n19 IBIAS.n6 20.3299
R5725 IBIAS.n17 IBIAS.n5 18.824
R5726 IBIAS.n15 IBIAS.n4 17.3181
R5727 IBIAS.n26 IBIAS.n2 16.3559
R5728 IBIAS.n13 IBIAS.n3 15.8123
R5729 IBIAS.n27 IBIAS.n1 12.7256
R5730 IBIAS.n11 IBIAS.n3 11.2946
R5731 IBIAS.n13 IBIAS.n4 9.78874
R5732 IBIAS.n1 IBIAS.n0 9.3005
R5733 IBIAS.n24 IBIAS.n23 9.3005
R5734 IBIAS.n22 IBIAS.n21 9.3005
R5735 IBIAS.n20 IBIAS.n19 9.3005
R5736 IBIAS.n18 IBIAS.n17 9.3005
R5737 IBIAS.n16 IBIAS.n15 9.3005
R5738 IBIAS.n14 IBIAS.n13 9.3005
R5739 IBIAS.n12 IBIAS.n11 9.3005
R5740 IBIAS.n15 IBIAS.n5 8.28285
R5741 IBIAS.n17 IBIAS.n6 6.77697
R5742 IBIAS.n19 IBIAS.n7 5.27109
R5743 IBIAS IBIAS.n28 5.23142
R5744 IBIAS.n21 IBIAS.n8 3.76521
R5745 IBIAS.n26 IBIAS.t2 2.48621
R5746 IBIAS.n26 IBIAS.t0 2.48621
R5747 IBIAS.n10 IBIAS.n2 2.36936
R5748 IBIAS.n25 IBIAS.n24 2.25932
R5749 IBIAS.n10 IBIAS.n9 0.320353
R5750 IBIAS.n28 IBIAS.n0 0.196152
R5751 IBIAS.n23 IBIAS.n0 0.196152
R5752 IBIAS.n23 IBIAS.n22 0.196152
R5753 IBIAS.n22 IBIAS.n20 0.196152
R5754 IBIAS.n20 IBIAS.n18 0.196152
R5755 IBIAS.n18 IBIAS.n16 0.196152
R5756 IBIAS.n16 IBIAS.n14 0.196152
R5757 IBIAS.n14 IBIAS.n12 0.196152
R5758 IBIAS.n12 IBIAS.n10 0.196152
C8 IBIAS VSS 2.04259f
C9 EN VSS 2.9958f
C10 VP VSS 5.00274f
C11 VN VSS 5.17776f
C12 VOUT VSS 20.55421f
C13 VDD VSS 14.42739f
C14 mim_cap_0.C1 VSS 33.98161f $ **FLOATING
C15 mim_cap_0.C1.t0 VSS 0.27321f $ **FLOATING
C16 mim_cap_0.C1.t1 VSS 28.5249f $ **FLOATING
C17 a_3758_2896.t6 VSS 0.03416f $ **FLOATING
C18 a_3758_2896.t3 VSS 0.03416f $ **FLOATING
C19 a_3758_2896.t4 VSS 0.03416f $ **FLOATING
C20 a_3758_2896.n0 VSS 0.11734f $ **FLOATING
C21 a_3758_2896.t0 VSS 0.03416f $ **FLOATING
C22 a_3758_2896.t10 VSS 0.03416f $ **FLOATING
C23 a_3758_2896.n1 VSS 0.10037f $ **FLOATING
C24 a_3758_2896.n2 VSS 0.75156f $ **FLOATING
C25 a_3758_2896.t9 VSS 0.03416f $ **FLOATING
C26 a_3758_2896.t8 VSS 0.03416f $ **FLOATING
C27 a_3758_2896.n3 VSS 0.10037f $ **FLOATING
C28 a_3758_2896.n4 VSS 0.39548f $ **FLOATING
C29 a_3758_2896.t2 VSS 0.03416f $ **FLOATING
C30 a_3758_2896.t1 VSS 0.03416f $ **FLOATING
C31 a_3758_2896.n5 VSS 0.10037f $ **FLOATING
C32 a_3758_2896.n6 VSS 0.39548f $ **FLOATING
C33 a_3758_2896.n7 VSS 0.01301f $ **FLOATING
C34 a_3758_2896.t13 VSS 0.12182f $ **FLOATING
C35 a_3758_2896.n9 VSS 0.01076f $ **FLOATING
C36 a_3758_2896.t12 VSS 0.79281f $ **FLOATING
C37 a_3758_2896.n16 VSS 1.50323f $ **FLOATING
C38 a_3758_2896.n17 VSS 0.21382f $ **FLOATING
C39 a_3758_2896.n19 VSS 0.01301f $ **FLOATING
C40 a_3758_2896.n21 VSS 0.01301f $ **FLOATING
C41 a_3758_2896.n23 VSS 0.01301f $ **FLOATING
C42 a_3758_2896.n25 VSS 0.01301f $ **FLOATING
C43 a_3758_2896.n27 VSS 0.01301f $ **FLOATING
C44 a_3758_2896.n29 VSS 0.01301f $ **FLOATING
C45 a_3758_2896.n30 VSS 0.01301f $ **FLOATING
C46 a_3758_2896.t14 VSS 0.07972f $ **FLOATING
C47 a_3758_2896.n33 VSS 0.17055f $ **FLOATING
C48 a_3758_2896.n35 VSS 0.36219f $ **FLOATING
C49 a_3758_2896.t5 VSS 0.03416f $ **FLOATING
C50 a_3758_2896.t7 VSS 0.03416f $ **FLOATING
C51 a_3758_2896.n36 VSS 0.10037f $ **FLOATING
C52 a_3758_2896.n37 VSS 0.64652f $ **FLOATING
C53 a_3758_2896.n38 VSS 0.33874f $ **FLOATING
C54 a_3758_2896.n39 VSS 0.10037f $ **FLOATING
C55 a_3758_2896.t11 VSS 0.03416f $ **FLOATING
C56 a_2479_9004.t3 VSS 1.50187f $ **FLOATING
C57 a_2479_9004.n0 VSS 2.87497f $ **FLOATING
C58 a_2479_9004.n5 VSS 0.01065f $ **FLOATING
C59 a_2479_9004.t18 VSS 0.15099f $ **FLOATING
C60 a_2479_9004.n9 VSS 0.40499f $ **FLOATING
C61 a_2479_9004.t12 VSS 0.02157f $ **FLOATING
C62 a_2479_9004.t10 VSS 0.02157f $ **FLOATING
C63 a_2479_9004.n10 VSS 0.04515f $ **FLOATING
C64 a_2479_9004.t8 VSS 0.02157f $ **FLOATING
C65 a_2479_9004.t6 VSS 0.02157f $ **FLOATING
C66 a_2479_9004.n11 VSS 0.04515f $ **FLOATING
C67 a_2479_9004.t23 VSS 0.09373f $ **FLOATING
C68 a_2479_9004.t7 VSS 0.09373f $ **FLOATING
C69 a_2479_9004.n13 VSS 0.23774f $ **FLOATING
C70 a_2479_9004.t24 VSS 0.09373f $ **FLOATING
C71 a_2479_9004.t5 VSS 0.09373f $ **FLOATING
C72 a_2479_9004.n14 VSS 0.24805f $ **FLOATING
C73 a_2479_9004.t11 VSS 0.09373f $ **FLOATING
C74 a_2479_9004.t21 VSS 0.09373f $ **FLOATING
C75 a_2479_9004.n15 VSS 0.24805f $ **FLOATING
C76 a_2479_9004.n16 VSS 0.23774f $ **FLOATING
C77 a_2479_9004.t9 VSS 0.09373f $ **FLOATING
C78 a_2479_9004.t22 VSS 0.09373f $ **FLOATING
C79 a_2479_9004.n17 VSS 0.94441f $ **FLOATING
C80 a_2479_9004.t16 VSS 0.15099f $ **FLOATING
C81 a_2479_9004.t15 VSS 0.15099f $ **FLOATING
C82 a_2479_9004.n18 VSS 0.83797f $ **FLOATING
C83 a_2479_9004.t20 VSS 0.15099f $ **FLOATING
C84 a_2479_9004.t19 VSS 0.15099f $ **FLOATING
C85 a_2479_9004.n19 VSS 0.6229f $ **FLOATING
C86 a_2479_9004.n20 VSS 3.08737f $ **FLOATING
C87 a_2479_9004.n21 VSS 1.8669f $ **FLOATING
C88 a_2479_9004.n22 VSS 0.02463f $ **FLOATING
C89 a_2479_9004.n23 VSS 0.01693f $ **FLOATING
C90 a_2479_9004.t17 VSS 0.15099f $ **FLOATING
C91 a_2479_9004.n24 VSS 0.02039f $ **FLOATING
C92 a_2479_9004.t2 VSS 0.07974f $ **FLOATING
C93 a_2479_9004.t0 VSS 1.50187f $ **FLOATING
C94 a_2479_9004.n31 VSS 2.87497f $ **FLOATING
C95 a_2479_9004.n32 VSS 0.40499f $ **FLOATING
C96 a_2479_9004.n33 VSS 0.01642f $ **FLOATING
C97 a_2479_9004.n34 VSS 0.02463f $ **FLOATING
C98 a_2479_9004.n36 VSS 0.02463f $ **FLOATING
C99 a_2479_9004.n38 VSS 0.02463f $ **FLOATING
C100 a_2479_9004.n40 VSS 0.02463f $ **FLOATING
C101 a_2479_9004.n42 VSS 0.02463f $ **FLOATING
C102 a_2479_9004.n44 VSS 0.02463f $ **FLOATING
C103 a_2479_9004.n45 VSS 0.02463f $ **FLOATING
C104 a_2479_9004.t1 VSS 0.15099f $ **FLOATING
C105 a_2479_9004.n48 VSS 0.32302f $ **FLOATING
C106 a_2479_9004.n49 VSS 0.01065f $ **FLOATING
C107 a_2479_9004.n50 VSS 0.37922f $ **FLOATING
C108 a_2479_9004.t14 VSS 0.15099f $ **FLOATING
C109 a_2479_9004.t13 VSS 0.15099f $ **FLOATING
C110 a_2479_9004.n51 VSS 0.60795f $ **FLOATING
C111 a_2479_9004.n52 VSS 1.42234f $ **FLOATING
C112 a_2479_9004.n53 VSS 0.3605f $ **FLOATING
C113 a_2479_9004.n54 VSS 0.19419f $ **FLOATING
C114 a_2479_9004.n55 VSS 0.01693f $ **FLOATING
C115 a_2479_9004.n56 VSS 0.02463f $ **FLOATING
C116 a_2479_9004.n58 VSS 0.02463f $ **FLOATING
C117 a_2479_9004.n60 VSS 0.02463f $ **FLOATING
C118 a_2479_9004.n62 VSS 0.02463f $ **FLOATING
C119 a_2479_9004.n64 VSS 0.02463f $ **FLOATING
C120 a_2479_9004.n66 VSS 0.02463f $ **FLOATING
C121 a_2479_9004.n68 VSS 0.02463f $ **FLOATING
C122 a_2479_9004.n69 VSS 0.02463f $ **FLOATING
C123 a_2479_9004.n70 VSS 0.01642f $ **FLOATING
C124 a_2479_9004.n71 VSS 0.02039f $ **FLOATING
C125 a_2479_9004.n72 VSS 0.32302f $ **FLOATING
C126 a_2479_9004.t4 VSS 0.23073f $ **FLOATING
C127 VN.t0 VSS 1.3922f $ **FLOATING
C128 VN.t1 VSS 1.38823f $ **FLOATING
C129 VN.n0 VSS 1.2253f $ **FLOATING
C130 VN.t4 VSS 1.38823f $ **FLOATING
C131 VN.n1 VSS 0.61184f $ **FLOATING
C132 VN.t5 VSS 1.38951f $ **FLOATING
C133 VN.n2 VSS 1.08963f $ **FLOATING
C134 VN.t7 VSS 1.38792f $ **FLOATING
C135 VN.t2 VSS 1.39115f $ **FLOATING
C136 VN.t6 VSS 1.38792f $ **FLOATING
C137 VN.n3 VSS 1.21058f $ **FLOATING
C138 VN.n4 VSS 0.57945f $ **FLOATING
C139 VN.t3 VSS 1.3877f $ **FLOATING
C140 VN.n5 VSS 0.60129f $ **FLOATING
C141 VN.n6 VSS 0.69029f $ **FLOATING
C142 a_2995_7336.t1 VSS 0.11279f $ **FLOATING
C143 a_2995_7336.t11 VSS 0.11279f $ **FLOATING
C144 a_2995_7336.t5 VSS 0.11279f $ **FLOATING
C145 a_2995_7336.n0 VSS 0.32272f $ **FLOATING
C146 a_2995_7336.t9 VSS 0.11279f $ **FLOATING
C147 a_2995_7336.t2 VSS 0.11279f $ **FLOATING
C148 a_2995_7336.n1 VSS 0.32268f $ **FLOATING
C149 a_2995_7336.t3 VSS 0.11279f $ **FLOATING
C150 a_2995_7336.t15 VSS 0.11279f $ **FLOATING
C151 a_2995_7336.n2 VSS 0.32272f $ **FLOATING
C152 a_2995_7336.n3 VSS 1.26812f $ **FLOATING
C153 a_2995_7336.n4 VSS 0.0184f $ **FLOATING
C154 a_2995_7336.n5 VSS 0.01264f $ **FLOATING
C155 a_2995_7336.t14 VSS 0.11279f $ **FLOATING
C156 a_2995_7336.n6 VSS 0.01523f $ **FLOATING
C157 a_2995_7336.t19 VSS 0.05957f $ **FLOATING
C158 a_2995_7336.t17 VSS 1.12173f $ **FLOATING
C159 a_2995_7336.n13 VSS 2.1269f $ **FLOATING
C160 a_2995_7336.n14 VSS 0.30254f $ **FLOATING
C161 a_2995_7336.n15 VSS 0.01227f $ **FLOATING
C162 a_2995_7336.n16 VSS 0.0184f $ **FLOATING
C163 a_2995_7336.n18 VSS 0.0184f $ **FLOATING
C164 a_2995_7336.n20 VSS 0.0184f $ **FLOATING
C165 a_2995_7336.n22 VSS 0.0184f $ **FLOATING
C166 a_2995_7336.n24 VSS 0.0184f $ **FLOATING
C167 a_2995_7336.n26 VSS 0.0184f $ **FLOATING
C168 a_2995_7336.n27 VSS 0.0184f $ **FLOATING
C169 a_2995_7336.t18 VSS 0.11279f $ **FLOATING
C170 a_2995_7336.n30 VSS 0.24131f $ **FLOATING
C171 a_2995_7336.n32 VSS 0.18922f $ **FLOATING
C172 a_2995_7336.t16 VSS 0.11279f $ **FLOATING
C173 a_2995_7336.t7 VSS 0.11279f $ **FLOATING
C174 a_2995_7336.n33 VSS 0.32268f $ **FLOATING
C175 a_2995_7336.t8 VSS 0.11279f $ **FLOATING
C176 a_2995_7336.t13 VSS 0.11279f $ **FLOATING
C177 a_2995_7336.n34 VSS 0.32272f $ **FLOATING
C178 a_2995_7336.t6 VSS 0.11279f $ **FLOATING
C179 a_2995_7336.t12 VSS 0.11279f $ **FLOATING
C180 a_2995_7336.n35 VSS 0.32268f $ **FLOATING
C181 a_2995_7336.t10 VSS 0.11279f $ **FLOATING
C182 a_2995_7336.t4 VSS 0.11279f $ **FLOATING
C183 a_2995_7336.n36 VSS 0.32272f $ **FLOATING
C184 a_2995_7336.n37 VSS 1.26812f $ **FLOATING
C185 a_2995_7336.n38 VSS 1.58502f $ **FLOATING
C186 a_2995_7336.n39 VSS 1.93909f $ **FLOATING
C187 a_2995_7336.n40 VSS 1.60505f $ **FLOATING
C188 a_2995_7336.n41 VSS 0.32272f $ **FLOATING
C189 a_2995_7336.t0 VSS 0.11279f $ **FLOATING
C190 VP.t7 VSS 1.39761f $ **FLOATING
C191 VP.t6 VSS 1.39363f $ **FLOATING
C192 VP.n0 VSS 1.23006f $ **FLOATING
C193 VP.t2 VSS 1.39363f $ **FLOATING
C194 VP.n1 VSS 0.61421f $ **FLOATING
C195 VP.t1 VSS 1.39491f $ **FLOATING
C196 VP.n2 VSS 1.09386f $ **FLOATING
C197 VP.t3 VSS 1.39656f $ **FLOATING
C198 VP.t5 VSS 1.39331f $ **FLOATING
C199 VP.n3 VSS 1.21529f $ **FLOATING
C200 VP.t4 VSS 1.39331f $ **FLOATING
C201 VP.n4 VSS 0.5817f $ **FLOATING
C202 VP.t0 VSS 1.39309f $ **FLOATING
C203 VP.n5 VSS 0.60363f $ **FLOATING
C204 VP.n6 VSS 0.6844f $ **FLOATING
C205 a_4920_2896.t10 VSS 0.02015f $ **FLOATING
C206 a_4920_2896.t16 VSS 0.02015f $ **FLOATING
C207 a_4920_2896.n0 VSS 0.04651f $ **FLOATING
C208 a_4920_2896.t4 VSS 0.02015f $ **FLOATING
C209 a_4920_2896.t11 VSS 0.02015f $ **FLOATING
C210 a_4920_2896.n1 VSS 0.04651f $ **FLOATING
C211 a_4920_2896.t20 VSS 0.02015f $ **FLOATING
C212 a_4920_2896.t3 VSS 0.02015f $ **FLOATING
C213 a_4920_2896.n2 VSS 0.04651f $ **FLOATING
C214 a_4920_2896.t22 VSS 0.02015f $ **FLOATING
C215 a_4920_2896.t21 VSS 0.02015f $ **FLOATING
C216 a_4920_2896.n3 VSS 0.04651f $ **FLOATING
C217 a_4920_2896.t14 VSS 0.02015f $ **FLOATING
C218 a_4920_2896.t9 VSS 0.02015f $ **FLOATING
C219 a_4920_2896.n4 VSS 0.05823f $ **FLOATING
C220 a_4920_2896.n5 VSS 0.44309f $ **FLOATING
C221 a_4920_2896.n6 VSS 0.18382f $ **FLOATING
C222 a_4920_2896.n7 VSS 0.18382f $ **FLOATING
C223 a_4920_2896.n8 VSS 0.18382f $ **FLOATING
C224 a_4920_2896.t8 VSS 0.02015f $ **FLOATING
C225 a_4920_2896.t1 VSS 0.02015f $ **FLOATING
C226 a_4920_2896.n9 VSS 0.04759f $ **FLOATING
C227 a_4920_2896.t18 VSS 0.02015f $ **FLOATING
C228 a_4920_2896.t2 VSS 0.02015f $ **FLOATING
C229 a_4920_2896.n10 VSS 0.04759f $ **FLOATING
C230 a_4920_2896.t13 VSS 0.02015f $ **FLOATING
C231 a_4920_2896.t19 VSS 0.02015f $ **FLOATING
C232 a_4920_2896.n11 VSS 0.04759f $ **FLOATING
C233 a_4920_2896.t5 VSS 0.02015f $ **FLOATING
C234 a_4920_2896.t12 VSS 0.02015f $ **FLOATING
C235 a_4920_2896.n12 VSS 0.04759f $ **FLOATING
C236 a_4920_2896.t7 VSS 0.02015f $ **FLOATING
C237 a_4920_2896.t6 VSS 0.02015f $ **FLOATING
C238 a_4920_2896.n13 VSS 0.04759f $ **FLOATING
C239 a_4920_2896.t0 VSS 0.02015f $ **FLOATING
C240 a_4920_2896.t17 VSS 0.02015f $ **FLOATING
C241 a_4920_2896.n14 VSS 0.05955f $ **FLOATING
C242 a_4920_2896.n15 VSS 0.4586f $ **FLOATING
C243 a_4920_2896.n16 VSS 0.1917f $ **FLOATING
C244 a_4920_2896.n17 VSS 0.1917f $ **FLOATING
C245 a_4920_2896.n18 VSS 0.1917f $ **FLOATING
C246 a_4920_2896.n19 VSS 0.37064f $ **FLOATING
C247 a_4920_2896.t26 VSS 0.07185f $ **FLOATING
C248 a_4920_2896.t25 VSS 0.46761f $ **FLOATING
C249 a_4920_2896.n30 VSS 0.88664f $ **FLOATING
C250 a_4920_2896.n44 VSS 0.12612f $ **FLOATING
C251 a_4920_2896.t24 VSS 0.04702f $ **FLOATING
C252 a_4920_2896.n46 VSS 0.10059f $ **FLOATING
C253 a_4920_2896.n48 VSS 0.0652f $ **FLOATING
C254 a_4920_2896.n49 VSS 0.31283f $ **FLOATING
C255 a_4920_2896.n50 VSS 0.23403f $ **FLOATING
C256 a_4920_2896.t15 VSS 0.02015f $ **FLOATING
C257 a_4920_2896.n51 VSS 0.04651f $ **FLOATING
C258 a_4920_2896.t23 VSS 0.02015f $ **FLOATING
C259 a_2080_2896.t2 VSS 0.02936f $ **FLOATING
C260 a_2080_2896.t3 VSS 0.01551f $ **FLOATING
C261 a_2080_2896.t1 VSS 0.29202f $ **FLOATING
C262 a_2080_2896.n9 VSS 0.5537f $ **FLOATING
C263 a_2080_2896.n10 VSS 0.07876f $ **FLOATING
C264 a_2080_2896.t22 VSS 0.21364f $ **FLOATING
C265 a_2080_2896.t30 VSS 0.21316f $ **FLOATING
C266 a_2080_2896.n24 VSS 0.22163f $ **FLOATING
C267 a_2080_2896.t9 VSS 0.21316f $ **FLOATING
C268 a_2080_2896.n25 VSS 0.08384f $ **FLOATING
C269 a_2080_2896.t10 VSS 0.21316f $ **FLOATING
C270 a_2080_2896.n26 VSS 0.08384f $ **FLOATING
C271 a_2080_2896.t11 VSS 0.21316f $ **FLOATING
C272 a_2080_2896.n27 VSS 0.08384f $ **FLOATING
C273 a_2080_2896.t40 VSS 0.21316f $ **FLOATING
C274 a_2080_2896.n28 VSS 0.08384f $ **FLOATING
C275 a_2080_2896.t39 VSS 0.21316f $ **FLOATING
C276 a_2080_2896.n29 VSS 0.08384f $ **FLOATING
C277 a_2080_2896.t28 VSS 0.21316f $ **FLOATING
C278 a_2080_2896.n30 VSS 0.08384f $ **FLOATING
C279 a_2080_2896.t29 VSS 0.21316f $ **FLOATING
C280 a_2080_2896.n31 VSS 0.08384f $ **FLOATING
C281 a_2080_2896.t18 VSS 0.21316f $ **FLOATING
C282 a_2080_2896.n32 VSS 0.08384f $ **FLOATING
C283 a_2080_2896.t8 VSS 0.21316f $ **FLOATING
C284 a_2080_2896.n33 VSS 0.08384f $ **FLOATING
C285 a_2080_2896.t21 VSS 0.21316f $ **FLOATING
C286 a_2080_2896.n34 VSS 0.11277f $ **FLOATING
C287 a_2080_2896.t35 VSS 0.21356f $ **FLOATING
C288 a_2080_2896.t43 VSS 0.21238f $ **FLOATING
C289 a_2080_2896.t27 VSS 0.21229f $ **FLOATING
C290 a_2080_2896.n35 VSS 0.1205f $ **FLOATING
C291 a_2080_2896.n36 VSS 0.13801f $ **FLOATING
C292 a_2080_2896.t15 VSS 0.21238f $ **FLOATING
C293 a_2080_2896.t38 VSS 0.21229f $ **FLOATING
C294 a_2080_2896.n37 VSS 0.1205f $ **FLOATING
C295 a_2080_2896.n38 VSS 0.02104f $ **FLOATING
C296 a_2080_2896.t32 VSS 0.21238f $ **FLOATING
C297 a_2080_2896.t16 VSS 0.21229f $ **FLOATING
C298 a_2080_2896.n39 VSS 0.1205f $ **FLOATING
C299 a_2080_2896.n40 VSS 0.02104f $ **FLOATING
C300 a_2080_2896.t33 VSS 0.21238f $ **FLOATING
C301 a_2080_2896.t17 VSS 0.21229f $ **FLOATING
C302 a_2080_2896.n41 VSS 0.1205f $ **FLOATING
C303 a_2080_2896.n42 VSS 0.02104f $ **FLOATING
C304 a_2080_2896.t34 VSS 0.21238f $ **FLOATING
C305 a_2080_2896.t19 VSS 0.21229f $ **FLOATING
C306 a_2080_2896.n43 VSS 0.1205f $ **FLOATING
C307 a_2080_2896.n44 VSS 0.02104f $ **FLOATING
C308 a_2080_2896.n45 VSS 0.02104f $ **FLOATING
C309 a_2080_2896.t23 VSS 0.21238f $ **FLOATING
C310 a_2080_2896.n46 VSS 0.01136f $ **FLOATING
C311 a_2080_2896.t25 VSS 0.21238f $ **FLOATING
C312 a_2080_2896.n47 VSS 0.07247f $ **FLOATING
C313 a_2080_2896.n48 VSS 0.04758f $ **FLOATING
C314 a_2080_2896.t6 VSS 0.16153f $ **FLOATING
C315 a_2080_2896.t7 VSS 0.01258f $ **FLOATING
C316 a_2080_2896.t5 VSS 0.01258f $ **FLOATING
C317 a_2080_2896.n68 VSS 0.02517f $ **FLOATING
C318 a_2080_2896.n71 VSS 0.11181f $ **FLOATING
C319 a_2080_2896.t4 VSS 0.16153f $ **FLOATING
C320 a_2080_2896.n72 VSS 0.04758f $ **FLOATING
C321 a_2080_2896.n73 VSS 0.07247f $ **FLOATING
C322 a_2080_2896.n74 VSS 0.02104f $ **FLOATING
C323 a_2080_2896.t12 VSS 0.21238f $ **FLOATING
C324 a_2080_2896.t36 VSS 0.21229f $ **FLOATING
C325 a_2080_2896.n75 VSS 0.1205f $ **FLOATING
C326 a_2080_2896.n76 VSS 0.02104f $ **FLOATING
C327 a_2080_2896.t13 VSS 0.21238f $ **FLOATING
C328 a_2080_2896.t37 VSS 0.21229f $ **FLOATING
C329 a_2080_2896.n77 VSS 0.1205f $ **FLOATING
C330 a_2080_2896.n78 VSS 0.02104f $ **FLOATING
C331 a_2080_2896.t41 VSS 0.21238f $ **FLOATING
C332 a_2080_2896.t24 VSS 0.21229f $ **FLOATING
C333 a_2080_2896.n79 VSS 0.1205f $ **FLOATING
C334 a_2080_2896.n80 VSS 0.02104f $ **FLOATING
C335 a_2080_2896.t31 VSS 0.21238f $ **FLOATING
C336 a_2080_2896.t14 VSS 0.21229f $ **FLOATING
C337 a_2080_2896.n81 VSS 0.1205f $ **FLOATING
C338 a_2080_2896.n82 VSS 0.02104f $ **FLOATING
C339 a_2080_2896.t42 VSS 0.21238f $ **FLOATING
C340 a_2080_2896.t26 VSS 0.21229f $ **FLOATING
C341 a_2080_2896.n83 VSS 0.1205f $ **FLOATING
C342 a_2080_2896.n84 VSS 0.02104f $ **FLOATING
C343 a_2080_2896.t20 VSS 0.21316f $ **FLOATING
C344 a_2080_2896.n85 VSS 0.16653f $ **FLOATING
C345 a_2080_2896.n86 VSS 0.2988f $ **FLOATING
C346 a_2080_2896.n87 VSS 0.17452f $ **FLOATING
C347 a_2080_2896.n91 VSS 0.06282f $ **FLOATING
C348 a_2080_2896.t0 VSS 0.02936f $ **FLOATING
C349 VDD.t18 VSS 0.03767f $ **FLOATING
C350 VDD.t64 VSS 0.01309f $ **FLOATING
C351 VDD.n0 VSS 0.0117f $ **FLOATING
C352 VDD.t16 VSS 0.03479f $ **FLOATING
C353 VDD.n1 VSS 0.20321f $ **FLOATING
C354 VDD.n2 VSS 0.01774f $ **FLOATING
C355 VDD.n3 VSS 0.18809f $ **FLOATING
C356 VDD.n4 VSS 0.01774f $ **FLOATING
C357 VDD.n5 VSS 0.12703f $ **FLOATING
C358 VDD.n6 VSS 0.01774f $ **FLOATING
C359 VDD.n7 VSS 0.12703f $ **FLOATING
C360 VDD.n8 VSS 0.01774f $ **FLOATING
C361 VDD.n9 VSS 0.16687f $ **FLOATING
C362 VDD.n10 VSS 0.05286f $ **FLOATING
C363 VDD.t12 VSS 0.01601f $ **FLOATING
C364 VDD.n11 VSS 0.02521f $ **FLOATING
C365 VDD.n12 VSS 0.02565f $ **FLOATING
C366 VDD.t24 VSS 0.03483f $ **FLOATING
C367 VDD.t35 VSS 0.06828f $ **FLOATING
C368 VDD.t36 VSS 0.03774f $ **FLOATING
C369 VDD.n13 VSS 0.04548f $ **FLOATING
C370 VDD.n14 VSS 0.01668f $ **FLOATING
C371 VDD.n15 VSS 0.02051f $ **FLOATING
C372 VDD.n16 VSS 0.07672f $ **FLOATING
C373 VDD.n17 VSS 0.04124f $ **FLOATING
C374 VDD.t10 VSS 0.06824f $ **FLOATING
C375 VDD.n18 VSS 0.02565f $ **FLOATING
C376 VDD.n19 VSS 0.04124f $ **FLOATING
C377 VDD.t46 VSS 0.06826f $ **FLOATING
C378 VDD.n20 VSS 0.0602f $ **FLOATING
C379 VDD.n21 VSS 0.01966f $ **FLOATING
C380 VDD.n22 VSS 0.02051f $ **FLOATING
C381 VDD.n23 VSS 0.01668f $ **FLOATING
C382 VDD.t48 VSS 0.01601f $ **FLOATING
C383 VDD.n24 VSS 0.0167f $ **FLOATING
C384 VDD.t26 VSS 0.01601f $ **FLOATING
C385 VDD.n25 VSS 0.0167f $ **FLOATING
C386 VDD.n26 VSS 0.10903f $ **FLOATING
C387 VDD.n27 VSS 0.01774f $ **FLOATING
C388 VDD.n28 VSS 0.24467f $ **FLOATING
C389 VDD.n29 VSS 0.05286f $ **FLOATING
C390 VDD.n30 VSS 0.02051f $ **FLOATING
C391 VDD.t9 VSS 0.02973f $ **FLOATING
C392 VDD.n31 VSS 0.07672f $ **FLOATING
C393 VDD.n32 VSS 0.02565f $ **FLOATING
C394 VDD.t49 VSS 0.03483f $ **FLOATING
C395 VDD.n33 VSS 0.01966f $ **FLOATING
C396 VDD.n34 VSS 0.0602f $ **FLOATING
C397 VDD.t27 VSS 0.06826f $ **FLOATING
C398 VDD.n35 VSS 0.02521f $ **FLOATING
C399 VDD.n36 VSS 0.04124f $ **FLOATING
C400 VDD.t30 VSS 0.06824f $ **FLOATING
C401 VDD.n37 VSS 0.02565f $ **FLOATING
C402 VDD.n38 VSS 0.04124f $ **FLOATING
C403 VDD.t6 VSS 0.06828f $ **FLOATING
C404 VDD.n39 VSS 0.04548f $ **FLOATING
C405 VDD.n40 VSS 0.02051f $ **FLOATING
C406 VDD.n41 VSS 0.01668f $ **FLOATING
C407 VDD.t32 VSS 0.01601f $ **FLOATING
C408 VDD.n42 VSS 0.01668f $ **FLOATING
C409 VDD.t29 VSS 0.01601f $ **FLOATING
C410 VDD.n43 VSS 0.0167f $ **FLOATING
C411 VDD.t50 VSS 0.01601f $ **FLOATING
C412 VDD.n44 VSS 0.0167f $ **FLOATING
C413 VDD.n45 VSS 0.08267f $ **FLOATING
C414 VDD.n46 VSS 0.07985f $ **FLOATING
C415 VDD.n52 VSS 0.52934f $ **FLOATING
C416 VDD.n65 VSS 0.01379f $ **FLOATING
C417 VDD.n68 VSS 0.01342f $ **FLOATING
C418 VDD.n71 VSS 0.36736f $ **FLOATING
C419 VDD.n73 VSS 0.01342f $ **FLOATING
C420 VDD.n76 VSS 0.37314f $ **FLOATING
C421 VDD.t31 VSS 0.19669f $ **FLOATING
C422 VDD.n80 VSS 0.37893f $ **FLOATING
C423 VDD.n84 VSS 0.38471f $ **FLOATING
C424 VDD.t14 VSS 0.19669f $ **FLOATING
C425 VDD.n88 VSS 0.3905f $ **FLOATING
C426 VDD.n92 VSS 0.39339f $ **FLOATING
C427 VDD.t55 VSS 0.19669f $ **FLOATING
C428 VDD.t2 VSS 0.19669f $ **FLOATING
C429 VDD.t0 VSS 0.19669f $ **FLOATING
C430 VDD.n99 VSS 0.3905f $ **FLOATING
C431 VDD.t25 VSS 0.19669f $ **FLOATING
C432 VDD.t47 VSS 0.19669f $ **FLOATING
C433 VDD.n106 VSS 0.37893f $ **FLOATING
C434 VDD.t11 VSS 0.19669f $ **FLOATING
C435 VDD.n111 VSS 0.01342f $ **FLOATING
C436 VDD.n112 VSS 0.01342f $ **FLOATING
C437 VDD.t17 VSS 0.19669f $ **FLOATING
C438 VDD.n113 VSS 0.36736f $ **FLOATING
C439 VDD.n114 VSS 0.01342f $ **FLOATING
C440 VDD.n116 VSS 0.52934f $ **FLOATING
C441 VDD.n117 VSS 0.67108f $ **FLOATING
C442 VDD.n125 VSS 0.01004f $ **FLOATING
C443 VDD.n136 VSS 0.01379f $ **FLOATING
C444 VDD.n137 VSS 0.01379f $ **FLOATING
C445 VDD.n157 VSS 0.01004f $ **FLOATING
C446 VDD.n158 VSS 0.01004f $ **FLOATING
C447 VDD.n159 VSS 0.01004f $ **FLOATING
C448 VDD.n180 VSS 0.01379f $ **FLOATING
C449 VDD.n181 VSS 0.01379f $ **FLOATING
C450 VDD.n182 VSS 0.01342f $ **FLOATING
C451 VDD.n185 VSS 0.22851f $ **FLOATING
C452 VDD.n191 VSS 0.37314f $ **FLOATING
C453 VDD.n192 VSS 0.22273f $ **FLOATING
C454 VDD.n198 VSS 0.21694f $ **FLOATING
C455 VDD.n204 VSS 0.38471f $ **FLOATING
C456 VDD.n205 VSS 0.21116f $ **FLOATING
C457 VDD.n211 VSS 0.20537f $ **FLOATING
C458 VDD.n217 VSS 0.19959f $ **FLOATING
C459 VDD.n223 VSS 0.19959f $ **FLOATING
C460 VDD.t4 VSS 0.19669f $ **FLOATING
C461 VDD.n229 VSS 0.20537f $ **FLOATING
C462 VDD.n235 VSS 0.21116f $ **FLOATING
C463 VDD.t28 VSS 0.19669f $ **FLOATING
C464 VDD.n241 VSS 0.21694f $ **FLOATING
C465 VDD.n247 VSS 0.22273f $ **FLOATING
C466 VDD.n255 VSS 0.01004f $ **FLOATING
C467 VDD.n256 VSS 0.01004f $ **FLOATING
C468 VDD.n257 VSS 0.01004f $ **FLOATING
C469 VDD.n258 VSS 0.01004f $ **FLOATING
C470 VDD.n281 VSS 0.01379f $ **FLOATING
C471 VDD.n282 VSS 0.01342f $ **FLOATING
C472 VDD.t7 VSS 0.19669f $ **FLOATING
C473 VDD.n285 VSS 0.22851f $ **FLOATING
C474 VDD.n288 VSS 0.01342f $ **FLOATING
C475 VDD.n296 VSS 0.01379f $ **FLOATING
C476 VDD.n297 VSS 0.01379f $ **FLOATING
C477 VDD.n299 VSS 0.67108f $ **FLOATING
C478 VDD.n304 VSS 0.0872f $ **FLOATING
C479 VDD.n305 VSS 0.07158f $ **FLOATING
C480 VDD.n306 VSS 0.05286f $ **FLOATING
C481 VDD.t23 VSS 0.01601f $ **FLOATING
C482 VDD.n307 VSS 0.01966f $ **FLOATING
C483 VDD.n308 VSS 0.07672f $ **FLOATING
C484 VDD.n309 VSS 0.04124f $ **FLOATING
C485 VDD.t44 VSS 0.06828f $ **FLOATING
C486 VDD.t45 VSS 0.03774f $ **FLOATING
C487 VDD.n310 VSS 0.01668f $ **FLOATING
C488 VDD.n311 VSS 0.02051f $ **FLOATING
C489 VDD.n312 VSS 0.04548f $ **FLOATING
C490 VDD.n313 VSS 0.02565f $ **FLOATING
C491 VDD.t22 VSS 0.06824f $ **FLOATING
C492 VDD.n314 VSS 0.02565f $ **FLOATING
C493 VDD.t33 VSS 0.03483f $ **FLOATING
C494 VDD.n315 VSS 0.0602f $ **FLOATING
C495 VDD.t51 VSS 0.06826f $ **FLOATING
C496 VDD.n316 VSS 0.04124f $ **FLOATING
C497 VDD.n317 VSS 0.02521f $ **FLOATING
C498 VDD.n318 VSS 0.02051f $ **FLOATING
C499 VDD.n319 VSS 0.01668f $ **FLOATING
C500 VDD.t52 VSS 0.01601f $ **FLOATING
C501 VDD.n320 VSS 0.0167f $ **FLOATING
C502 VDD.t34 VSS 0.01601f $ **FLOATING
C503 VDD.n321 VSS 0.0167f $ **FLOATING
C504 VDD.n322 VSS 0.1092f $ **FLOATING
C505 VDD.n323 VSS 0.01774f $ **FLOATING
C506 VDD.n324 VSS 0.24543f $ **FLOATING
C507 VDD.n325 VSS 0.05286f $ **FLOATING
C508 VDD.n326 VSS 0.02051f $ **FLOATING
C509 VDD.n327 VSS 0.04548f $ **FLOATING
C510 VDD.n328 VSS 0.02521f $ **FLOATING
C511 VDD.t21 VSS 0.02973f $ **FLOATING
C512 VDD.n329 VSS 0.04124f $ **FLOATING
C513 VDD.t13 VSS 0.03483f $ **FLOATING
C514 VDD.t37 VSS 0.06826f $ **FLOATING
C515 VDD.n330 VSS 0.0602f $ **FLOATING
C516 VDD.n331 VSS 0.01966f $ **FLOATING
C517 VDD.n332 VSS 0.02565f $ **FLOATING
C518 VDD.t42 VSS 0.06824f $ **FLOATING
C519 VDD.n333 VSS 0.02565f $ **FLOATING
C520 VDD.t19 VSS 0.06828f $ **FLOATING
C521 VDD.n334 VSS 0.04124f $ **FLOATING
C522 VDD.n335 VSS 0.07672f $ **FLOATING
C523 VDD.n336 VSS 0.02051f $ **FLOATING
C524 VDD.n337 VSS 0.01668f $ **FLOATING
C525 VDD.t43 VSS 0.01601f $ **FLOATING
C526 VDD.n338 VSS 0.01668f $ **FLOATING
C527 VDD.t38 VSS 0.01601f $ **FLOATING
C528 VDD.n339 VSS 0.0167f $ **FLOATING
C529 VDD.t15 VSS 0.01601f $ **FLOATING
C530 VDD.n340 VSS 0.0167f $ **FLOATING
C531 VDD.n341 VSS 0.08267f $ **FLOATING
C532 VDD.n342 VSS 0.10025f $ **FLOATING
C533 VDD.n343 VSS 0.01833f $ **FLOATING
C534 VDD.n344 VSS 0.01774f $ **FLOATING
C535 VDD.n345 VSS 0.3241f $ **FLOATING
C536 VDD.n346 VSS 0.01774f $ **FLOATING
C537 VDD.n347 VSS 0.12703f $ **FLOATING
C538 VDD.n348 VSS 0.01774f $ **FLOATING
C539 VDD.n349 VSS 0.12703f $ **FLOATING
C540 VDD.t41 VSS 0.02967f $ **FLOATING
C541 VDD.n350 VSS 0.0167f $ **FLOATING
C542 VDD.n351 VSS 0.11338f $ **FLOATING
C543 VDD.t39 VSS 0.03479f $ **FLOATING
C544 VDD.n352 VSS 0.07466f $ **FLOATING
C545 VDD.n353 VSS 0.10377f $ **FLOATING
C546 VDD.n354 VSS 0.41757f $ **FLOATING
C547 VDD.n355 VSS 0.27238f $ **FLOATING
C548 VDD.n356 VSS 0.17089f $ **FLOATING
C549 VOUT.n0 VSS 0.01561f $ **FLOATING
C550 VOUT.n1 VSS 0.01513f $ **FLOATING
C551 VOUT.n2 VSS 0.2765f $ **FLOATING
C552 VOUT.n3 VSS 0.01513f $ **FLOATING
C553 VOUT.n4 VSS 0.11605f $ **FLOATING
C554 VOUT.n5 VSS 0.01513f $ **FLOATING
C555 VOUT.n6 VSS 0.11605f $ **FLOATING
C556 VOUT.n7 VSS 0.03194f $ **FLOATING
C557 VOUT.n8 VSS 0.03838f $ **FLOATING
C558 VOUT.t26 VSS 0.05763f $ **FLOATING
C559 VOUT.t28 VSS 0.02509f $ **FLOATING
C560 VOUT.n9 VSS 0.01408f $ **FLOATING
C561 VOUT.t23 VSS 0.01351f $ **FLOATING
C562 VOUT.n10 VSS 0.01408f $ **FLOATING
C563 VOUT.n11 VSS 0.01731f $ **FLOATING
C564 VOUT.n12 VSS 0.06898f $ **FLOATING
C565 VOUT.n13 VSS 0.0566f $ **FLOATING
C566 VOUT.t22 VSS 0.05761f $ **FLOATING
C567 VOUT.n14 VSS 0.02164f $ **FLOATING
C568 VOUT.n15 VSS 0.04613f $ **FLOATING
C569 VOUT.n16 VSS 0.10296f $ **FLOATING
C570 VOUT.t0 VSS 0.04729f $ **FLOATING
C571 VOUT.t31 VSS 0.02497f $ **FLOATING
C572 VOUT.t29 VSS 0.47028f $ **FLOATING
C573 VOUT.n26 VSS 0.89169f $ **FLOATING
C574 VOUT.n27 VSS 0.12684f $ **FLOATING
C575 VOUT.t30 VSS 0.04729f $ **FLOATING
C576 VOUT.n43 VSS 0.10117f $ **FLOATING
C577 VOUT.n45 VSS 0.44202f $ **FLOATING
C578 VOUT.n46 VSS 0.66282f $ **FLOATING
C579 VOUT.t19 VSS 67.909f $ **FLOATING
C580 VOUT.n47 VSS 0.26662f $ **FLOATING
C581 VOUT.n48 VSS 0.02041f $ **FLOATING
C582 VOUT.n49 VSS 0.06898f $ **FLOATING
C583 VOUT.t21 VSS 0.03185f $ **FLOATING
C584 VOUT.t24 VSS 0.05761f $ **FLOATING
C585 VOUT.n50 VSS 0.0566f $ **FLOATING
C586 VOUT.t20 VSS 0.05763f $ **FLOATING
C587 VOUT.n51 VSS 0.03838f $ **FLOATING
C588 VOUT.n52 VSS 0.01731f $ **FLOATING
C589 VOUT.n53 VSS 0.01408f $ **FLOATING
C590 VOUT.t25 VSS 0.01351f $ **FLOATING
C591 VOUT.n54 VSS 0.01408f $ **FLOATING
C592 VOUT.n55 VSS 0.0334f $ **FLOATING
C593 VOUT.n56 VSS 0.06133f $ **FLOATING
C594 VOUT.n57 VSS 0.01513f $ **FLOATING
C595 VOUT.n58 VSS 0.18517f $ **FLOATING
C596 VOUT.n59 VSS 0.01513f $ **FLOATING
C597 VOUT.n60 VSS 0.11605f $ **FLOATING
C598 VOUT.n61 VSS 0.01513f $ **FLOATING
C599 VOUT.n62 VSS 0.11605f $ **FLOATING
C600 VOUT.n63 VSS 0.01513f $ **FLOATING
C601 VOUT.n64 VSS 0.16056f $ **FLOATING
C602 VOUT.n65 VSS 0.27398f $ **FLOATING
C603 VOUT.n66 VSS 0.3823f $ **FLOATING
C604 a_2479_7336.t11 VSS 0.11568f $ **FLOATING
C605 a_2479_7336.t13 VSS 0.01653f $ **FLOATING
C606 a_2479_7336.t14 VSS 0.01653f $ **FLOATING
C607 a_2479_7336.n0 VSS 0.03485f $ **FLOATING
C608 a_2479_7336.t31 VSS 0.07191f $ **FLOATING
C609 a_2479_7336.t22 VSS 0.07182f $ **FLOATING
C610 a_2479_7336.n1 VSS 0.13333f $ **FLOATING
C611 a_2479_7336.t24 VSS 0.07182f $ **FLOATING
C612 a_2479_7336.n2 VSS 0.06199f $ **FLOATING
C613 a_2479_7336.n3 VSS 0.16118f $ **FLOATING
C614 a_2479_7336.t27 VSS 0.07182f $ **FLOATING
C615 a_2479_7336.n4 VSS 0.06199f $ **FLOATING
C616 a_2479_7336.t33 VSS 0.07182f $ **FLOATING
C617 a_2479_7336.n5 VSS 0.07104f $ **FLOATING
C618 a_2479_7336.t18 VSS 0.07182f $ **FLOATING
C619 a_2479_7336.n6 VSS 0.07104f $ **FLOATING
C620 a_2479_7336.t29 VSS 0.07182f $ **FLOATING
C621 a_2479_7336.n7 VSS 0.07104f $ **FLOATING
C622 a_2479_7336.t21 VSS 0.07182f $ **FLOATING
C623 a_2479_7336.n8 VSS 0.07104f $ **FLOATING
C624 a_2479_7336.t34 VSS 0.07182f $ **FLOATING
C625 a_2479_7336.n9 VSS 0.12436f $ **FLOATING
C626 a_2479_7336.t15 VSS 0.01653f $ **FLOATING
C627 a_2479_7336.t3 VSS 0.01653f $ **FLOATING
C628 a_2479_7336.n10 VSS 0.03485f $ **FLOATING
C629 a_2479_7336.t19 VSS 0.07191f $ **FLOATING
C630 a_2479_7336.t28 VSS 0.07182f $ **FLOATING
C631 a_2479_7336.n11 VSS 0.13333f $ **FLOATING
C632 a_2479_7336.t35 VSS 0.07182f $ **FLOATING
C633 a_2479_7336.n12 VSS 0.06199f $ **FLOATING
C634 a_2479_7336.n13 VSS 0.16118f $ **FLOATING
C635 a_2479_7336.t32 VSS 0.07182f $ **FLOATING
C636 a_2479_7336.n14 VSS 0.06199f $ **FLOATING
C637 a_2479_7336.t26 VSS 0.07182f $ **FLOATING
C638 a_2479_7336.n15 VSS 0.07104f $ **FLOATING
C639 a_2479_7336.t23 VSS 0.07182f $ **FLOATING
C640 a_2479_7336.n16 VSS 0.07104f $ **FLOATING
C641 a_2479_7336.t20 VSS 0.07182f $ **FLOATING
C642 a_2479_7336.n17 VSS 0.07104f $ **FLOATING
C643 a_2479_7336.t30 VSS 0.07182f $ **FLOATING
C644 a_2479_7336.n18 VSS 0.07104f $ **FLOATING
C645 a_2479_7336.t25 VSS 0.07182f $ **FLOATING
C646 a_2479_7336.n19 VSS 0.12097f $ **FLOATING
C647 a_2479_7336.t17 VSS 0.71057f $ **FLOATING
C648 a_2479_7336.n20 VSS 4.9407f $ **FLOATING
C649 a_2479_7336.n21 VSS 2.25646f $ **FLOATING
C650 a_2479_7336.t2 VSS 0.11568f $ **FLOATING
C651 a_2479_7336.t1 VSS 0.11568f $ **FLOATING
C652 a_2479_7336.n22 VSS 0.47727f $ **FLOATING
C653 a_2479_7336.n23 VSS 1.44242f $ **FLOATING
C654 a_2479_7336.n24 VSS 0.01887f $ **FLOATING
C655 a_2479_7336.n25 VSS 0.01297f $ **FLOATING
C656 a_2479_7336.t8 VSS 0.17677f $ **FLOATING
C657 a_2479_7336.n33 VSS 0.01258f $ **FLOATING
C658 a_2479_7336.t7 VSS 1.15067f $ **FLOATING
C659 a_2479_7336.n34 VSS 2.20269f $ **FLOATING
C660 a_2479_7336.n36 VSS 0.01887f $ **FLOATING
C661 a_2479_7336.n38 VSS 0.01887f $ **FLOATING
C662 a_2479_7336.n40 VSS 0.01887f $ **FLOATING
C663 a_2479_7336.n42 VSS 0.01887f $ **FLOATING
C664 a_2479_7336.n44 VSS 0.01887f $ **FLOATING
C665 a_2479_7336.n46 VSS 0.01887f $ **FLOATING
C666 a_2479_7336.n47 VSS 0.01887f $ **FLOATING
C667 a_2479_7336.n48 VSS 0.31029f $ **FLOATING
C668 a_2479_7336.n49 VSS 0.01562f $ **FLOATING
C669 a_2479_7336.t12 VSS 0.11568f $ **FLOATING
C670 a_2479_7336.n50 VSS 0.24749f $ **FLOATING
C671 a_2479_7336.n52 VSS 0.29048f $ **FLOATING
C672 a_2479_7336.t9 VSS 0.11568f $ **FLOATING
C673 a_2479_7336.t16 VSS 0.11568f $ **FLOATING
C674 a_2479_7336.n53 VSS 0.46576f $ **FLOATING
C675 a_2479_7336.n54 VSS 1.08983f $ **FLOATING
C676 a_2479_7336.n55 VSS 0.01887f $ **FLOATING
C677 a_2479_7336.n56 VSS 0.01297f $ **FLOATING
C678 a_2479_7336.t10 VSS 0.11568f $ **FLOATING
C679 a_2479_7336.n64 VSS 0.01258f $ **FLOATING
C680 a_2479_7336.t6 VSS 0.06109f $ **FLOATING
C681 a_2479_7336.t4 VSS 1.15067f $ **FLOATING
C682 a_2479_7336.n65 VSS 2.20269f $ **FLOATING
C683 a_2479_7336.n67 VSS 0.01887f $ **FLOATING
C684 a_2479_7336.n69 VSS 0.01887f $ **FLOATING
C685 a_2479_7336.n71 VSS 0.01887f $ **FLOATING
C686 a_2479_7336.n73 VSS 0.01887f $ **FLOATING
C687 a_2479_7336.n75 VSS 0.01887f $ **FLOATING
C688 a_2479_7336.n77 VSS 0.01887f $ **FLOATING
C689 a_2479_7336.n78 VSS 0.01887f $ **FLOATING
C690 a_2479_7336.n79 VSS 0.31029f $ **FLOATING
C691 a_2479_7336.n80 VSS 0.01562f $ **FLOATING
C692 a_2479_7336.t5 VSS 0.11568f $ **FLOATING
C693 a_2479_7336.n81 VSS 0.24749f $ **FLOATING
C694 a_2479_7336.n83 VSS 0.14878f $ **FLOATING
C695 a_2479_7336.n84 VSS 1.03586f $ **FLOATING
C696 a_2479_7336.n85 VSS 1.60671f $ **FLOATING
C697 a_2479_7336.n86 VSS 0.47725f $ **FLOATING
C698 a_2479_7336.t0 VSS 0.11568f $ **FLOATING
.ends
