VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_lochidev_two_stage_opamp
  CLASS BLOCK ;
  FOREIGN tt_um_lochidev_two_stage_opamp ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 7.000000 ;
    ANTENNADIFFAREA 4.060000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 226.000000 ;
    ANTENNADIFFAREA 122.163795 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 85.599998 ;
    ANTENNADIFFAREA 8.120000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNAGATEAREA 85.599998 ;
    ANTENNADIFFAREA 8.120000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 85.599998 ;
    ANTENNADIFFAREA 8.120000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 7.200000 ;
    ANTENNADIFFAREA 16.445799 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 32.730 67.470 52.450 67.900 ;
        RECT 32.730 65.360 33.160 67.470 ;
        RECT 52.020 65.360 52.450 67.470 ;
        RECT 32.730 64.930 52.450 65.360 ;
        RECT 11.755 53.230 26.225 61.360 ;
      LAYER nwell ;
        RECT 32.185 54.135 42.135 64.615 ;
      LAYER pwell ;
        RECT 11.755 52.150 12.185 53.230 ;
        RECT 25.795 52.150 26.225 53.230 ;
        RECT 11.755 44.890 26.225 52.150 ;
        RECT 11.755 43.810 12.185 44.890 ;
        RECT 25.795 43.810 26.225 44.890 ;
        RECT 11.755 36.550 26.225 43.810 ;
        RECT 11.755 35.470 12.185 36.550 ;
        RECT 25.795 35.470 26.225 36.550 ;
        RECT 11.755 27.340 26.225 35.470 ;
        RECT 9.760 13.480 26.820 22.480 ;
        RECT 28.895 22.295 51.105 26.425 ;
        RECT 28.895 20.795 29.325 22.295 ;
        RECT 50.675 20.795 51.105 22.295 ;
        RECT 28.895 17.535 51.105 20.795 ;
        RECT 28.895 16.035 29.325 17.535 ;
        RECT 50.675 16.035 51.105 17.535 ;
        RECT 28.895 11.905 51.105 16.035 ;
      LAYER li1 ;
        RECT 32.860 67.600 52.320 67.770 ;
        RECT 32.860 65.230 33.030 67.600 ;
        RECT 33.510 65.710 35.670 67.120 ;
        RECT 49.510 65.710 51.670 67.120 ;
        RECT 52.150 65.230 52.320 67.600 ;
        RECT 32.860 65.060 52.320 65.230 ;
        RECT 32.365 64.265 41.955 64.435 ;
        RECT 11.885 61.060 26.095 61.230 ;
        RECT 11.885 27.640 12.055 61.060 ;
        RECT 12.685 60.550 13.685 60.720 ;
        RECT 13.975 60.550 14.975 60.720 ;
        RECT 15.265 60.550 16.265 60.720 ;
        RECT 16.555 60.550 17.555 60.720 ;
        RECT 17.845 60.550 18.845 60.720 ;
        RECT 19.135 60.550 20.135 60.720 ;
        RECT 20.425 60.550 21.425 60.720 ;
        RECT 21.715 60.550 22.715 60.720 ;
        RECT 23.005 60.550 24.005 60.720 ;
        RECT 24.295 60.550 25.295 60.720 ;
        RECT 12.455 53.340 12.625 60.380 ;
        RECT 13.745 53.340 13.915 60.380 ;
        RECT 15.035 53.340 15.205 60.380 ;
        RECT 16.325 53.340 16.495 60.380 ;
        RECT 17.615 53.340 17.785 60.380 ;
        RECT 18.905 53.340 19.075 60.380 ;
        RECT 20.195 53.340 20.365 60.380 ;
        RECT 21.485 53.340 21.655 60.380 ;
        RECT 22.775 53.340 22.945 60.380 ;
        RECT 24.065 53.340 24.235 60.380 ;
        RECT 25.355 53.340 25.525 60.380 ;
        RECT 12.685 52.210 13.685 52.380 ;
        RECT 13.975 52.210 14.975 52.380 ;
        RECT 15.265 52.210 16.265 52.380 ;
        RECT 16.555 52.210 17.555 52.380 ;
        RECT 17.845 52.210 18.845 52.380 ;
        RECT 19.135 52.210 20.135 52.380 ;
        RECT 20.425 52.210 21.425 52.380 ;
        RECT 21.715 52.210 22.715 52.380 ;
        RECT 23.005 52.210 24.005 52.380 ;
        RECT 24.295 52.210 25.295 52.380 ;
        RECT 12.455 45.000 12.625 52.040 ;
        RECT 13.745 45.000 13.915 52.040 ;
        RECT 15.035 45.000 15.205 52.040 ;
        RECT 16.325 45.000 16.495 52.040 ;
        RECT 17.615 45.000 17.785 52.040 ;
        RECT 18.905 45.000 19.075 52.040 ;
        RECT 20.195 45.000 20.365 52.040 ;
        RECT 21.485 45.000 21.655 52.040 ;
        RECT 22.775 45.000 22.945 52.040 ;
        RECT 24.065 45.000 24.235 52.040 ;
        RECT 25.355 45.000 25.525 52.040 ;
        RECT 12.685 44.660 13.685 44.830 ;
        RECT 13.975 44.660 14.975 44.830 ;
        RECT 15.265 44.660 16.265 44.830 ;
        RECT 16.555 44.660 17.555 44.830 ;
        RECT 17.845 44.660 18.845 44.830 ;
        RECT 19.135 44.660 20.135 44.830 ;
        RECT 20.425 44.660 21.425 44.830 ;
        RECT 21.715 44.660 22.715 44.830 ;
        RECT 23.005 44.660 24.005 44.830 ;
        RECT 24.295 44.660 25.295 44.830 ;
        RECT 12.685 43.870 13.685 44.040 ;
        RECT 13.975 43.870 14.975 44.040 ;
        RECT 15.265 43.870 16.265 44.040 ;
        RECT 16.555 43.870 17.555 44.040 ;
        RECT 17.845 43.870 18.845 44.040 ;
        RECT 19.135 43.870 20.135 44.040 ;
        RECT 20.425 43.870 21.425 44.040 ;
        RECT 21.715 43.870 22.715 44.040 ;
        RECT 23.005 43.870 24.005 44.040 ;
        RECT 24.295 43.870 25.295 44.040 ;
        RECT 12.455 36.660 12.625 43.700 ;
        RECT 13.745 36.660 13.915 43.700 ;
        RECT 15.035 36.660 15.205 43.700 ;
        RECT 16.325 36.660 16.495 43.700 ;
        RECT 17.615 36.660 17.785 43.700 ;
        RECT 18.905 36.660 19.075 43.700 ;
        RECT 20.195 36.660 20.365 43.700 ;
        RECT 21.485 36.660 21.655 43.700 ;
        RECT 22.775 36.660 22.945 43.700 ;
        RECT 24.065 36.660 24.235 43.700 ;
        RECT 25.355 36.660 25.525 43.700 ;
        RECT 12.685 36.320 13.685 36.490 ;
        RECT 13.975 36.320 14.975 36.490 ;
        RECT 15.265 36.320 16.265 36.490 ;
        RECT 16.555 36.320 17.555 36.490 ;
        RECT 17.845 36.320 18.845 36.490 ;
        RECT 19.135 36.320 20.135 36.490 ;
        RECT 20.425 36.320 21.425 36.490 ;
        RECT 21.715 36.320 22.715 36.490 ;
        RECT 23.005 36.320 24.005 36.490 ;
        RECT 24.295 36.320 25.295 36.490 ;
        RECT 12.455 28.320 12.625 35.360 ;
        RECT 13.745 28.320 13.915 35.360 ;
        RECT 15.035 28.320 15.205 35.360 ;
        RECT 16.325 28.320 16.495 35.360 ;
        RECT 17.615 28.320 17.785 35.360 ;
        RECT 18.905 28.320 19.075 35.360 ;
        RECT 20.195 28.320 20.365 35.360 ;
        RECT 21.485 28.320 21.655 35.360 ;
        RECT 22.775 28.320 22.945 35.360 ;
        RECT 24.065 28.320 24.235 35.360 ;
        RECT 25.355 28.320 25.525 35.360 ;
        RECT 12.685 27.980 13.685 28.150 ;
        RECT 13.975 27.980 14.975 28.150 ;
        RECT 15.265 27.980 16.265 28.150 ;
        RECT 16.555 27.980 17.555 28.150 ;
        RECT 17.845 27.980 18.845 28.150 ;
        RECT 19.135 27.980 20.135 28.150 ;
        RECT 20.425 27.980 21.425 28.150 ;
        RECT 21.715 27.980 22.715 28.150 ;
        RECT 23.005 27.980 24.005 28.150 ;
        RECT 24.295 27.980 25.295 28.150 ;
        RECT 25.925 27.640 26.095 61.060 ;
        RECT 32.365 54.485 32.535 64.265 ;
        RECT 33.165 63.755 33.565 63.925 ;
        RECT 33.855 63.755 34.255 63.925 ;
        RECT 40.755 63.755 41.155 63.925 ;
        RECT 32.935 62.500 33.105 63.540 ;
        RECT 33.625 62.500 33.795 63.540 ;
        RECT 34.315 62.500 34.485 63.540 ;
        RECT 35.005 62.500 35.175 63.540 ;
        RECT 35.695 62.500 35.865 63.540 ;
        RECT 36.385 62.500 36.555 63.540 ;
        RECT 37.075 62.500 37.245 63.540 ;
        RECT 37.765 62.500 37.935 63.540 ;
        RECT 38.455 62.500 38.625 63.540 ;
        RECT 39.145 62.500 39.315 63.540 ;
        RECT 39.835 62.500 40.005 63.540 ;
        RECT 40.525 62.500 40.695 63.540 ;
        RECT 41.215 62.500 41.385 63.540 ;
        RECT 33.165 62.115 33.565 62.285 ;
        RECT 33.855 62.115 34.255 62.285 ;
        RECT 34.545 62.115 34.945 62.285 ;
        RECT 35.235 62.115 35.635 62.285 ;
        RECT 35.925 62.115 36.325 62.285 ;
        RECT 36.615 62.115 37.015 62.285 ;
        RECT 37.305 62.115 37.705 62.285 ;
        RECT 37.995 62.115 38.395 62.285 ;
        RECT 38.685 62.115 39.085 62.285 ;
        RECT 39.375 62.115 39.775 62.285 ;
        RECT 40.065 62.115 40.465 62.285 ;
        RECT 33.165 61.325 33.565 61.495 ;
        RECT 33.855 61.325 34.255 61.495 ;
        RECT 34.545 61.325 34.945 61.495 ;
        RECT 39.375 61.325 39.775 61.495 ;
        RECT 40.065 61.325 40.465 61.495 ;
        RECT 40.755 61.325 41.155 61.495 ;
        RECT 32.935 60.070 33.105 61.110 ;
        RECT 33.625 60.070 33.795 61.110 ;
        RECT 34.315 60.070 34.485 61.110 ;
        RECT 35.005 60.070 35.175 61.110 ;
        RECT 35.695 60.070 35.865 61.110 ;
        RECT 36.385 60.070 36.555 61.110 ;
        RECT 37.075 60.070 37.245 61.110 ;
        RECT 37.765 60.070 37.935 61.110 ;
        RECT 38.455 60.070 38.625 61.110 ;
        RECT 39.145 60.070 39.315 61.110 ;
        RECT 39.835 60.070 40.005 61.110 ;
        RECT 40.525 60.070 40.695 61.110 ;
        RECT 41.215 60.070 41.385 61.110 ;
        RECT 33.165 59.685 33.565 59.855 ;
        RECT 33.855 59.685 34.255 59.855 ;
        RECT 34.545 59.685 34.945 59.855 ;
        RECT 35.235 59.685 35.635 59.855 ;
        RECT 35.925 59.685 36.325 59.855 ;
        RECT 36.615 59.685 37.015 59.855 ;
        RECT 37.305 59.685 37.705 59.855 ;
        RECT 37.995 59.685 38.395 59.855 ;
        RECT 38.685 59.685 39.085 59.855 ;
        RECT 39.375 59.685 39.775 59.855 ;
        RECT 40.065 59.685 40.465 59.855 ;
        RECT 40.755 59.685 41.155 59.855 ;
        RECT 33.165 58.895 33.565 59.065 ;
        RECT 33.855 58.895 34.255 59.065 ;
        RECT 34.545 58.895 34.945 59.065 ;
        RECT 35.235 58.895 35.635 59.065 ;
        RECT 35.925 58.895 36.325 59.065 ;
        RECT 36.615 58.895 37.015 59.065 ;
        RECT 37.305 58.895 37.705 59.065 ;
        RECT 37.995 58.895 38.395 59.065 ;
        RECT 38.685 58.895 39.085 59.065 ;
        RECT 39.375 58.895 39.775 59.065 ;
        RECT 40.065 58.895 40.465 59.065 ;
        RECT 40.755 58.895 41.155 59.065 ;
        RECT 32.935 57.640 33.105 58.680 ;
        RECT 33.625 57.640 33.795 58.680 ;
        RECT 34.315 57.640 34.485 58.680 ;
        RECT 35.005 57.640 35.175 58.680 ;
        RECT 35.695 57.640 35.865 58.680 ;
        RECT 36.385 57.640 36.555 58.680 ;
        RECT 37.075 57.640 37.245 58.680 ;
        RECT 37.765 57.640 37.935 58.680 ;
        RECT 38.455 57.640 38.625 58.680 ;
        RECT 39.145 57.640 39.315 58.680 ;
        RECT 39.835 57.640 40.005 58.680 ;
        RECT 40.525 57.640 40.695 58.680 ;
        RECT 41.215 57.640 41.385 58.680 ;
        RECT 33.165 57.255 33.565 57.425 ;
        RECT 33.855 57.255 34.255 57.425 ;
        RECT 34.545 57.255 34.945 57.425 ;
        RECT 39.375 57.255 39.775 57.425 ;
        RECT 40.065 57.255 40.465 57.425 ;
        RECT 40.755 57.255 41.155 57.425 ;
        RECT 33.855 56.465 34.255 56.635 ;
        RECT 34.545 56.465 34.945 56.635 ;
        RECT 35.235 56.465 35.635 56.635 ;
        RECT 35.925 56.465 36.325 56.635 ;
        RECT 36.615 56.465 37.015 56.635 ;
        RECT 37.305 56.465 37.705 56.635 ;
        RECT 37.995 56.465 38.395 56.635 ;
        RECT 38.685 56.465 39.085 56.635 ;
        RECT 39.375 56.465 39.775 56.635 ;
        RECT 40.065 56.465 40.465 56.635 ;
        RECT 40.755 56.465 41.155 56.635 ;
        RECT 32.935 55.210 33.105 56.250 ;
        RECT 33.625 55.210 33.795 56.250 ;
        RECT 34.315 55.210 34.485 56.250 ;
        RECT 35.005 55.210 35.175 56.250 ;
        RECT 35.695 55.210 35.865 56.250 ;
        RECT 36.385 55.210 36.555 56.250 ;
        RECT 37.075 55.210 37.245 56.250 ;
        RECT 37.765 55.210 37.935 56.250 ;
        RECT 38.455 55.210 38.625 56.250 ;
        RECT 39.145 55.210 39.315 56.250 ;
        RECT 39.835 55.210 40.005 56.250 ;
        RECT 40.525 55.210 40.695 56.250 ;
        RECT 41.215 55.210 41.385 56.250 ;
        RECT 33.165 54.825 33.565 54.995 ;
        RECT 40.065 54.825 40.465 54.995 ;
        RECT 40.755 54.825 41.155 54.995 ;
        RECT 41.785 54.485 41.955 64.265 ;
        RECT 32.365 54.315 41.955 54.485 ;
        RECT 11.885 27.470 26.095 27.640 ;
        RECT 29.025 26.125 50.975 26.295 ;
        RECT 9.890 22.180 15.070 22.350 ;
        RECT 9.890 13.780 10.060 22.180 ;
        RECT 10.690 21.670 11.690 21.840 ;
        RECT 11.980 21.670 12.980 21.840 ;
        RECT 13.270 21.670 14.270 21.840 ;
        RECT 10.460 14.460 10.630 21.500 ;
        RECT 11.750 14.460 11.920 21.500 ;
        RECT 13.040 14.460 13.210 21.500 ;
        RECT 14.330 14.460 14.500 21.500 ;
        RECT 10.690 14.120 11.690 14.290 ;
        RECT 11.980 14.120 12.980 14.290 ;
        RECT 13.270 14.120 14.270 14.290 ;
        RECT 14.900 13.780 15.070 22.180 ;
        RECT 9.890 13.610 15.070 13.780 ;
        RECT 15.700 22.180 20.880 22.350 ;
        RECT 15.700 13.780 15.870 22.180 ;
        RECT 16.500 21.670 17.500 21.840 ;
        RECT 17.790 21.670 18.790 21.840 ;
        RECT 19.080 21.670 20.080 21.840 ;
        RECT 16.270 14.460 16.440 21.500 ;
        RECT 17.560 14.460 17.730 21.500 ;
        RECT 18.850 14.460 19.020 21.500 ;
        RECT 20.140 14.460 20.310 21.500 ;
        RECT 16.500 14.120 17.500 14.290 ;
        RECT 17.790 14.120 18.790 14.290 ;
        RECT 19.080 14.120 20.080 14.290 ;
        RECT 20.710 13.780 20.880 22.180 ;
        RECT 15.700 13.610 20.880 13.780 ;
        RECT 21.510 22.180 26.690 22.350 ;
        RECT 21.510 13.780 21.680 22.180 ;
        RECT 22.310 21.670 23.310 21.840 ;
        RECT 23.600 21.670 24.600 21.840 ;
        RECT 24.890 21.670 25.890 21.840 ;
        RECT 22.080 14.460 22.250 21.500 ;
        RECT 23.370 14.460 23.540 21.500 ;
        RECT 24.660 14.460 24.830 21.500 ;
        RECT 25.950 14.460 26.120 21.500 ;
        RECT 22.310 14.120 23.310 14.290 ;
        RECT 23.600 14.120 24.600 14.290 ;
        RECT 24.890 14.120 25.890 14.290 ;
        RECT 26.520 13.780 26.690 22.180 ;
        RECT 21.510 13.610 26.690 13.780 ;
        RECT 29.025 12.205 29.195 26.125 ;
        RECT 29.825 25.615 30.825 25.785 ;
        RECT 31.115 25.615 32.115 25.785 ;
        RECT 32.405 25.615 33.405 25.785 ;
        RECT 33.695 25.615 34.695 25.785 ;
        RECT 34.985 25.615 35.985 25.785 ;
        RECT 36.275 25.615 37.275 25.785 ;
        RECT 37.565 25.615 38.565 25.785 ;
        RECT 38.855 25.615 39.855 25.785 ;
        RECT 40.145 25.615 41.145 25.785 ;
        RECT 41.435 25.615 42.435 25.785 ;
        RECT 42.725 25.615 43.725 25.785 ;
        RECT 44.015 25.615 45.015 25.785 ;
        RECT 45.305 25.615 46.305 25.785 ;
        RECT 46.595 25.615 47.595 25.785 ;
        RECT 47.885 25.615 48.885 25.785 ;
        RECT 49.175 25.615 50.175 25.785 ;
        RECT 29.595 22.405 29.765 25.445 ;
        RECT 30.885 22.405 31.055 25.445 ;
        RECT 32.175 22.405 32.345 25.445 ;
        RECT 33.465 22.405 33.635 25.445 ;
        RECT 34.755 22.405 34.925 25.445 ;
        RECT 36.045 22.405 36.215 25.445 ;
        RECT 37.335 22.405 37.505 25.445 ;
        RECT 38.625 22.405 38.795 25.445 ;
        RECT 39.915 22.405 40.085 25.445 ;
        RECT 41.205 22.405 41.375 25.445 ;
        RECT 42.495 22.405 42.665 25.445 ;
        RECT 43.785 22.405 43.955 25.445 ;
        RECT 45.075 22.405 45.245 25.445 ;
        RECT 46.365 22.405 46.535 25.445 ;
        RECT 47.655 22.405 47.825 25.445 ;
        RECT 48.945 22.405 49.115 25.445 ;
        RECT 50.235 22.405 50.405 25.445 ;
        RECT 29.825 22.065 30.825 22.235 ;
        RECT 31.115 22.065 32.115 22.235 ;
        RECT 32.405 22.065 33.405 22.235 ;
        RECT 33.695 22.065 34.695 22.235 ;
        RECT 34.985 22.065 35.985 22.235 ;
        RECT 36.275 22.065 37.275 22.235 ;
        RECT 37.565 22.065 38.565 22.235 ;
        RECT 38.855 22.065 39.855 22.235 ;
        RECT 40.145 22.065 41.145 22.235 ;
        RECT 41.435 22.065 42.435 22.235 ;
        RECT 42.725 22.065 43.725 22.235 ;
        RECT 44.015 22.065 45.015 22.235 ;
        RECT 45.305 22.065 46.305 22.235 ;
        RECT 46.595 22.065 47.595 22.235 ;
        RECT 47.885 22.065 48.885 22.235 ;
        RECT 49.175 22.065 50.175 22.235 ;
        RECT 29.825 20.855 30.825 21.025 ;
        RECT 31.115 20.855 32.115 21.025 ;
        RECT 32.405 20.855 33.405 21.025 ;
        RECT 33.695 20.855 34.695 21.025 ;
        RECT 34.985 20.855 35.985 21.025 ;
        RECT 36.275 20.855 37.275 21.025 ;
        RECT 37.565 20.855 38.565 21.025 ;
        RECT 38.855 20.855 39.855 21.025 ;
        RECT 40.145 20.855 41.145 21.025 ;
        RECT 41.435 20.855 42.435 21.025 ;
        RECT 42.725 20.855 43.725 21.025 ;
        RECT 44.015 20.855 45.015 21.025 ;
        RECT 45.305 20.855 46.305 21.025 ;
        RECT 46.595 20.855 47.595 21.025 ;
        RECT 47.885 20.855 48.885 21.025 ;
        RECT 49.175 20.855 50.175 21.025 ;
        RECT 29.595 17.645 29.765 20.685 ;
        RECT 30.885 17.645 31.055 20.685 ;
        RECT 32.175 17.645 32.345 20.685 ;
        RECT 33.465 17.645 33.635 20.685 ;
        RECT 34.755 17.645 34.925 20.685 ;
        RECT 36.045 17.645 36.215 20.685 ;
        RECT 37.335 17.645 37.505 20.685 ;
        RECT 38.625 17.645 38.795 20.685 ;
        RECT 39.915 17.645 40.085 20.685 ;
        RECT 41.205 17.645 41.375 20.685 ;
        RECT 42.495 17.645 42.665 20.685 ;
        RECT 43.785 17.645 43.955 20.685 ;
        RECT 45.075 17.645 45.245 20.685 ;
        RECT 46.365 17.645 46.535 20.685 ;
        RECT 47.655 17.645 47.825 20.685 ;
        RECT 48.945 17.645 49.115 20.685 ;
        RECT 50.235 17.645 50.405 20.685 ;
        RECT 29.825 17.305 30.825 17.475 ;
        RECT 31.115 17.305 32.115 17.475 ;
        RECT 32.405 17.305 33.405 17.475 ;
        RECT 33.695 17.305 34.695 17.475 ;
        RECT 34.985 17.305 35.985 17.475 ;
        RECT 36.275 17.305 37.275 17.475 ;
        RECT 37.565 17.305 38.565 17.475 ;
        RECT 38.855 17.305 39.855 17.475 ;
        RECT 40.145 17.305 41.145 17.475 ;
        RECT 41.435 17.305 42.435 17.475 ;
        RECT 42.725 17.305 43.725 17.475 ;
        RECT 44.015 17.305 45.015 17.475 ;
        RECT 45.305 17.305 46.305 17.475 ;
        RECT 46.595 17.305 47.595 17.475 ;
        RECT 47.885 17.305 48.885 17.475 ;
        RECT 49.175 17.305 50.175 17.475 ;
        RECT 29.825 16.095 30.825 16.265 ;
        RECT 31.115 16.095 32.115 16.265 ;
        RECT 32.405 16.095 33.405 16.265 ;
        RECT 33.695 16.095 34.695 16.265 ;
        RECT 34.985 16.095 35.985 16.265 ;
        RECT 36.275 16.095 37.275 16.265 ;
        RECT 37.565 16.095 38.565 16.265 ;
        RECT 38.855 16.095 39.855 16.265 ;
        RECT 40.145 16.095 41.145 16.265 ;
        RECT 41.435 16.095 42.435 16.265 ;
        RECT 42.725 16.095 43.725 16.265 ;
        RECT 44.015 16.095 45.015 16.265 ;
        RECT 45.305 16.095 46.305 16.265 ;
        RECT 46.595 16.095 47.595 16.265 ;
        RECT 47.885 16.095 48.885 16.265 ;
        RECT 49.175 16.095 50.175 16.265 ;
        RECT 29.595 12.885 29.765 15.925 ;
        RECT 30.885 12.885 31.055 15.925 ;
        RECT 32.175 12.885 32.345 15.925 ;
        RECT 33.465 12.885 33.635 15.925 ;
        RECT 34.755 12.885 34.925 15.925 ;
        RECT 36.045 12.885 36.215 15.925 ;
        RECT 37.335 12.885 37.505 15.925 ;
        RECT 38.625 12.885 38.795 15.925 ;
        RECT 39.915 12.885 40.085 15.925 ;
        RECT 41.205 12.885 41.375 15.925 ;
        RECT 42.495 12.885 42.665 15.925 ;
        RECT 43.785 12.885 43.955 15.925 ;
        RECT 45.075 12.885 45.245 15.925 ;
        RECT 46.365 12.885 46.535 15.925 ;
        RECT 47.655 12.885 47.825 15.925 ;
        RECT 48.945 12.885 49.115 15.925 ;
        RECT 50.235 12.885 50.405 15.925 ;
        RECT 29.825 12.545 30.825 12.715 ;
        RECT 31.115 12.545 32.115 12.715 ;
        RECT 32.405 12.545 33.405 12.715 ;
        RECT 33.695 12.545 34.695 12.715 ;
        RECT 34.985 12.545 35.985 12.715 ;
        RECT 36.275 12.545 37.275 12.715 ;
        RECT 37.565 12.545 38.565 12.715 ;
        RECT 38.855 12.545 39.855 12.715 ;
        RECT 40.145 12.545 41.145 12.715 ;
        RECT 41.435 12.545 42.435 12.715 ;
        RECT 42.725 12.545 43.725 12.715 ;
        RECT 44.015 12.545 45.015 12.715 ;
        RECT 45.305 12.545 46.305 12.715 ;
        RECT 46.595 12.545 47.595 12.715 ;
        RECT 47.885 12.545 48.885 12.715 ;
        RECT 49.175 12.545 50.175 12.715 ;
        RECT 50.805 12.205 50.975 26.125 ;
        RECT 29.025 12.035 50.975 12.205 ;
      LAYER met1 ;
        RECT 7.660 68.260 33.085 69.165 ;
        RECT 7.660 19.955 9.310 68.260 ;
        RECT 30.500 63.775 31.280 66.890 ;
        RECT 32.805 66.025 33.085 68.260 ;
        RECT 33.540 65.615 35.645 67.070 ;
        RECT 49.535 65.760 53.820 67.070 ;
        RECT 33.540 64.935 43.460 65.615 ;
        RECT 33.970 64.515 34.830 64.795 ;
        RECT 35.350 64.515 36.210 64.795 ;
        RECT 36.730 64.515 37.590 64.795 ;
        RECT 38.110 64.515 38.970 64.795 ;
        RECT 39.490 64.515 40.350 64.795 ;
        RECT 34.285 63.955 34.515 64.515 ;
        RECT 34.660 64.095 35.520 64.375 ;
        RECT 33.185 63.725 34.515 63.955 ;
        RECT 31.935 61.945 32.660 63.575 ;
        RECT 32.905 62.925 33.135 63.520 ;
        RECT 33.595 62.925 33.825 63.725 ;
        RECT 34.285 62.925 34.515 63.725 ;
        RECT 32.905 62.755 34.515 62.925 ;
        RECT 32.905 62.520 33.135 62.755 ;
        RECT 33.595 62.315 33.825 62.755 ;
        RECT 34.285 62.520 34.515 62.755 ;
        RECT 34.975 62.520 35.205 64.095 ;
        RECT 35.665 62.520 35.895 64.515 ;
        RECT 36.040 64.095 36.900 64.375 ;
        RECT 36.355 62.520 36.585 64.095 ;
        RECT 37.045 62.520 37.275 64.515 ;
        RECT 37.420 64.095 38.280 64.375 ;
        RECT 37.735 62.520 37.965 64.095 ;
        RECT 38.425 62.520 38.655 64.515 ;
        RECT 38.800 64.095 39.660 64.375 ;
        RECT 39.115 62.520 39.345 64.095 ;
        RECT 39.805 62.520 40.035 64.515 ;
        RECT 40.180 64.095 41.040 64.375 ;
        RECT 40.495 63.955 40.725 64.095 ;
        RECT 40.495 63.755 41.135 63.955 ;
        RECT 40.495 63.520 41.185 63.755 ;
        RECT 40.495 63.115 41.415 63.520 ;
        RECT 40.495 62.520 40.725 63.115 ;
        RECT 41.185 62.520 41.415 63.115 ;
        RECT 42.860 62.315 43.460 64.935 ;
        RECT 33.185 62.085 34.235 62.315 ;
        RECT 34.565 62.085 43.460 62.315 ;
        RECT 31.935 61.665 32.880 61.945 ;
        RECT 35.350 61.665 36.210 61.945 ;
        RECT 13.540 61.285 14.120 61.355 ;
        RECT 18.700 61.285 19.280 61.355 ;
        RECT 23.860 61.285 24.440 61.355 ;
        RECT 12.470 61.005 15.190 61.285 ;
        RECT 17.630 61.005 20.350 61.285 ;
        RECT 22.790 61.005 25.510 61.285 ;
        RECT 13.540 60.935 14.120 61.005 ;
        RECT 18.700 60.935 19.280 61.005 ;
        RECT 23.860 60.935 24.440 61.005 ;
        RECT 13.665 60.750 13.995 60.935 ;
        RECT 18.825 60.750 19.155 60.935 ;
        RECT 23.985 60.750 24.315 60.935 ;
        RECT 12.705 60.520 25.275 60.750 ;
        RECT 12.425 60.185 12.655 60.360 ;
        RECT 13.715 60.185 13.945 60.520 ;
        RECT 15.005 60.185 15.235 60.360 ;
        RECT 16.295 60.185 16.525 60.360 ;
        RECT 17.585 60.185 17.815 60.360 ;
        RECT 18.875 60.185 19.105 60.520 ;
        RECT 20.165 60.185 20.395 60.360 ;
        RECT 21.455 60.185 21.685 60.360 ;
        RECT 22.745 60.185 22.975 60.360 ;
        RECT 24.035 60.185 24.265 60.520 ;
        RECT 25.325 60.185 25.555 60.360 ;
        RECT 12.425 60.015 25.555 60.185 ;
        RECT 31.935 60.035 32.660 61.665 ;
        RECT 33.185 61.295 34.925 61.525 ;
        RECT 32.905 60.855 33.135 61.090 ;
        RECT 33.595 60.855 33.825 61.295 ;
        RECT 34.285 60.855 34.515 61.295 ;
        RECT 34.975 60.855 35.205 61.090 ;
        RECT 35.665 60.855 35.895 61.665 ;
        RECT 32.905 60.685 35.895 60.855 ;
        RECT 32.905 60.090 33.135 60.685 ;
        RECT 12.425 53.360 12.655 60.015 ;
        RECT 12.795 53.390 13.575 53.670 ;
        RECT 13.160 52.830 13.390 53.390 ;
        RECT 13.715 53.360 13.945 60.015 ;
        RECT 15.005 53.360 15.235 60.015 ;
        RECT 15.375 53.810 16.155 54.090 ;
        RECT 14.085 53.185 14.865 53.250 ;
        RECT 14.085 53.035 15.435 53.185 ;
        RECT 14.085 52.970 14.865 53.035 ;
        RECT 9.475 52.050 11.340 52.830 ;
        RECT 11.480 44.490 11.760 52.830 ;
        RECT 13.160 52.600 13.945 52.830 ;
        RECT 12.705 52.180 13.575 52.410 ;
        RECT 12.425 48.605 12.655 52.020 ;
        RECT 13.090 48.605 13.280 52.180 ;
        RECT 13.715 48.605 13.945 52.600 ;
        RECT 14.085 52.550 14.865 52.830 ;
        RECT 14.380 52.410 14.570 52.550 ;
        RECT 15.285 52.410 15.435 53.035 ;
        RECT 15.740 52.830 15.970 53.810 ;
        RECT 16.295 53.360 16.525 60.015 ;
        RECT 17.585 53.360 17.815 60.015 ;
        RECT 18.875 53.360 19.105 60.015 ;
        RECT 19.245 53.390 20.025 53.670 ;
        RECT 16.665 52.970 17.445 53.250 ;
        RECT 15.740 52.600 16.525 52.830 ;
        RECT 14.085 52.180 14.955 52.410 ;
        RECT 15.285 52.180 16.155 52.410 ;
        RECT 12.425 48.435 13.945 48.605 ;
        RECT 12.425 45.020 12.655 48.435 ;
        RECT 13.090 44.860 13.280 48.435 ;
        RECT 13.715 45.020 13.945 48.435 ;
        RECT 12.705 44.630 13.665 44.860 ;
        RECT 13.995 44.630 14.865 44.860 ;
        RECT 15.005 44.490 15.235 52.020 ;
        RECT 16.295 45.020 16.525 52.600 ;
        RECT 16.960 52.410 17.150 52.970 ;
        RECT 19.430 52.830 19.660 53.390 ;
        RECT 20.165 53.360 20.395 60.015 ;
        RECT 21.455 53.360 21.685 60.015 ;
        RECT 21.825 53.810 22.605 54.090 ;
        RECT 20.535 52.970 21.315 53.250 ;
        RECT 17.290 52.550 18.080 52.830 ;
        RECT 17.865 52.410 18.080 52.550 ;
        RECT 18.875 52.600 19.660 52.830 ;
        RECT 16.665 52.180 17.535 52.410 ;
        RECT 17.865 52.180 18.735 52.410 ;
        RECT 15.375 44.630 16.245 44.860 ;
        RECT 16.575 44.630 17.445 44.860 ;
        RECT 17.585 44.490 17.815 52.020 ;
        RECT 18.875 45.020 19.105 52.600 ;
        RECT 19.900 52.550 20.690 52.830 ;
        RECT 19.900 52.410 20.115 52.550 ;
        RECT 20.830 52.410 21.020 52.970 ;
        RECT 22.010 52.830 22.240 53.810 ;
        RECT 22.745 53.360 22.975 60.015 ;
        RECT 24.035 53.360 24.265 60.015 ;
        RECT 24.405 53.390 25.185 53.670 ;
        RECT 23.115 53.185 23.895 53.250 ;
        RECT 21.455 52.600 22.240 52.830 ;
        RECT 22.545 53.035 23.895 53.185 ;
        RECT 19.245 52.180 20.115 52.410 ;
        RECT 20.445 52.180 21.315 52.410 ;
        RECT 17.955 44.630 18.825 44.860 ;
        RECT 19.155 44.630 20.025 44.860 ;
        RECT 20.165 44.490 20.395 52.020 ;
        RECT 21.455 45.020 21.685 52.600 ;
        RECT 22.545 52.410 22.695 53.035 ;
        RECT 23.115 52.970 23.895 53.035 ;
        RECT 24.590 52.830 24.820 53.390 ;
        RECT 25.325 53.360 25.555 60.015 ;
        RECT 27.060 59.515 27.340 59.900 ;
        RECT 33.595 59.885 33.825 60.685 ;
        RECT 34.285 59.885 34.515 60.685 ;
        RECT 34.975 60.090 35.205 60.685 ;
        RECT 35.665 60.090 35.895 60.685 ;
        RECT 36.355 60.090 36.585 62.085 ;
        RECT 36.730 61.665 37.590 61.945 ;
        RECT 38.110 61.665 38.970 61.945 ;
        RECT 37.045 60.090 37.275 61.665 ;
        RECT 37.735 59.885 37.965 61.090 ;
        RECT 38.425 60.855 38.655 61.665 ;
        RECT 39.395 61.295 41.135 61.525 ;
        RECT 39.115 60.855 39.345 61.090 ;
        RECT 39.805 60.855 40.035 61.295 ;
        RECT 40.495 60.855 40.725 61.295 ;
        RECT 41.185 60.855 41.415 61.090 ;
        RECT 38.425 60.685 41.415 60.855 ;
        RECT 41.660 60.765 42.385 61.945 ;
        RECT 38.425 60.090 38.655 60.685 ;
        RECT 39.115 60.090 39.345 60.685 ;
        RECT 39.805 59.885 40.035 60.685 ;
        RECT 40.495 59.885 40.725 60.685 ;
        RECT 41.185 60.090 41.415 60.685 ;
        RECT 33.185 59.655 35.615 59.885 ;
        RECT 35.945 59.515 38.375 59.885 ;
        RECT 38.705 59.655 41.135 59.885 ;
        RECT 27.060 59.235 42.605 59.515 ;
        RECT 27.060 58.770 27.340 59.235 ;
        RECT 33.185 58.865 35.615 59.095 ;
        RECT 35.945 58.865 38.375 59.235 ;
        RECT 38.705 58.865 41.135 59.095 ;
        RECT 32.905 58.065 33.135 58.660 ;
        RECT 33.595 58.065 33.825 58.865 ;
        RECT 34.285 58.065 34.515 58.865 ;
        RECT 34.975 58.065 35.205 58.660 ;
        RECT 35.665 58.065 35.895 58.660 ;
        RECT 32.905 57.895 35.895 58.065 ;
        RECT 32.905 57.660 33.135 57.895 ;
        RECT 33.595 57.455 33.825 57.895 ;
        RECT 34.285 57.455 34.515 57.895 ;
        RECT 34.975 57.660 35.205 57.895 ;
        RECT 33.185 57.225 34.925 57.455 ;
        RECT 35.665 57.085 35.895 57.895 ;
        RECT 36.355 57.660 36.585 58.865 ;
        RECT 37.045 57.085 37.275 58.660 ;
        RECT 35.350 56.805 36.210 57.085 ;
        RECT 36.730 56.805 37.590 57.085 ;
        RECT 37.735 56.665 37.965 58.660 ;
        RECT 38.425 58.065 38.655 58.660 ;
        RECT 39.115 58.065 39.345 58.660 ;
        RECT 39.805 58.065 40.035 58.865 ;
        RECT 40.495 58.065 40.725 58.865 ;
        RECT 41.185 58.065 41.415 58.660 ;
        RECT 38.425 57.895 41.415 58.065 ;
        RECT 38.425 57.085 38.655 57.895 ;
        RECT 39.115 57.660 39.345 57.895 ;
        RECT 39.805 57.455 40.035 57.895 ;
        RECT 40.495 57.455 40.725 57.895 ;
        RECT 41.185 57.660 41.415 57.895 ;
        RECT 39.395 57.225 41.135 57.455 ;
        RECT 38.110 56.805 38.970 57.085 ;
        RECT 31.270 56.435 39.755 56.665 ;
        RECT 40.085 56.435 41.135 56.665 ;
        RECT 26.640 55.825 26.920 56.255 ;
        RECT 31.270 55.825 31.930 56.435 ;
        RECT 26.640 55.655 31.930 55.825 ;
        RECT 26.640 55.125 26.920 55.655 ;
        RECT 27.785 53.420 30.715 53.700 ;
        RECT 23.115 52.550 23.895 52.830 ;
        RECT 24.035 52.600 24.820 52.830 ;
        RECT 23.410 52.410 23.600 52.550 ;
        RECT 21.825 52.180 22.695 52.410 ;
        RECT 23.025 52.180 23.895 52.410 ;
        RECT 20.535 44.630 21.405 44.860 ;
        RECT 21.735 44.630 22.605 44.860 ;
        RECT 22.745 44.490 22.975 52.020 ;
        RECT 24.035 48.605 24.265 52.600 ;
        RECT 24.405 52.180 25.275 52.410 ;
        RECT 24.700 48.605 24.890 52.180 ;
        RECT 25.325 48.605 25.555 52.020 ;
        RECT 24.035 48.435 25.555 48.605 ;
        RECT 24.035 45.020 24.265 48.435 ;
        RECT 24.700 44.860 24.890 48.435 ;
        RECT 25.325 45.020 25.555 48.435 ;
        RECT 23.115 44.630 23.985 44.860 ;
        RECT 24.315 44.630 25.275 44.860 ;
        RECT 26.220 44.490 26.500 53.200 ;
        RECT 11.480 44.210 26.500 44.490 ;
        RECT 11.480 27.105 11.760 44.210 ;
        RECT 12.705 43.840 13.665 44.070 ;
        RECT 13.995 43.840 14.865 44.070 ;
        RECT 12.425 40.265 12.655 43.680 ;
        RECT 13.090 40.265 13.280 43.840 ;
        RECT 13.715 40.265 13.945 43.680 ;
        RECT 12.425 40.095 13.945 40.265 ;
        RECT 12.425 36.680 12.655 40.095 ;
        RECT 13.090 36.520 13.280 40.095 ;
        RECT 12.705 36.290 13.575 36.520 ;
        RECT 13.715 36.100 13.945 40.095 ;
        RECT 15.005 36.680 15.235 44.210 ;
        RECT 15.375 43.840 16.245 44.070 ;
        RECT 16.575 43.840 17.445 44.070 ;
        RECT 14.085 36.290 14.955 36.520 ;
        RECT 15.285 36.290 16.155 36.520 ;
        RECT 14.380 36.150 14.570 36.290 ;
        RECT 13.160 35.870 13.945 36.100 ;
        RECT 14.085 35.870 14.865 36.150 ;
        RECT 12.425 28.685 12.655 35.340 ;
        RECT 13.160 35.310 13.390 35.870 ;
        RECT 14.085 35.665 14.865 35.730 ;
        RECT 15.285 35.665 15.435 36.290 ;
        RECT 16.295 36.100 16.525 43.680 ;
        RECT 17.585 36.680 17.815 44.210 ;
        RECT 17.955 43.840 18.825 44.070 ;
        RECT 19.155 43.840 20.025 44.070 ;
        RECT 16.665 36.290 17.535 36.520 ;
        RECT 17.865 36.290 18.735 36.520 ;
        RECT 14.085 35.515 15.435 35.665 ;
        RECT 15.740 35.870 16.525 36.100 ;
        RECT 14.085 35.450 14.865 35.515 ;
        RECT 12.795 35.030 13.575 35.310 ;
        RECT 13.715 28.685 13.945 35.340 ;
        RECT 15.005 28.685 15.235 35.340 ;
        RECT 15.740 34.890 15.970 35.870 ;
        RECT 16.960 35.730 17.150 36.290 ;
        RECT 17.865 36.150 18.080 36.290 ;
        RECT 17.290 35.870 18.080 36.150 ;
        RECT 18.875 36.100 19.105 43.680 ;
        RECT 20.165 36.680 20.395 44.210 ;
        RECT 20.535 43.840 21.405 44.070 ;
        RECT 21.735 43.840 22.605 44.070 ;
        RECT 19.245 36.290 20.115 36.520 ;
        RECT 20.445 36.290 21.315 36.520 ;
        RECT 18.320 35.870 19.105 36.100 ;
        RECT 19.900 36.150 20.115 36.290 ;
        RECT 19.900 35.870 20.690 36.150 ;
        RECT 16.665 35.450 17.445 35.730 ;
        RECT 15.375 34.610 16.155 34.890 ;
        RECT 16.295 28.685 16.525 35.340 ;
        RECT 17.585 28.685 17.815 35.340 ;
        RECT 18.320 35.310 18.550 35.870 ;
        RECT 20.830 35.730 21.020 36.290 ;
        RECT 21.455 36.100 21.685 43.680 ;
        RECT 22.745 36.680 22.975 44.210 ;
        RECT 23.115 43.840 23.985 44.070 ;
        RECT 24.315 43.840 25.275 44.070 ;
        RECT 24.035 40.265 24.265 43.680 ;
        RECT 24.700 40.265 24.890 43.840 ;
        RECT 25.325 40.265 25.555 43.680 ;
        RECT 24.035 40.095 25.555 40.265 ;
        RECT 21.825 36.290 22.695 36.520 ;
        RECT 23.025 36.290 23.895 36.520 ;
        RECT 21.455 35.870 22.240 36.100 ;
        RECT 20.535 35.450 21.315 35.730 ;
        RECT 17.955 35.030 18.735 35.310 ;
        RECT 18.875 28.685 19.105 35.340 ;
        RECT 20.165 28.685 20.395 35.340 ;
        RECT 21.455 28.685 21.685 35.340 ;
        RECT 22.010 34.890 22.240 35.870 ;
        RECT 22.545 35.665 22.695 36.290 ;
        RECT 23.410 36.150 23.600 36.290 ;
        RECT 23.115 35.870 23.895 36.150 ;
        RECT 24.035 36.100 24.265 40.095 ;
        RECT 24.700 36.520 24.890 40.095 ;
        RECT 25.325 36.680 25.555 40.095 ;
        RECT 24.405 36.290 25.275 36.520 ;
        RECT 24.035 35.870 24.820 36.100 ;
        RECT 23.115 35.665 23.895 35.730 ;
        RECT 22.545 35.515 23.895 35.665 ;
        RECT 23.115 35.450 23.895 35.515 ;
        RECT 21.825 34.610 22.605 34.890 ;
        RECT 22.745 28.685 22.975 35.340 ;
        RECT 24.035 28.685 24.265 35.340 ;
        RECT 24.590 35.310 24.820 35.870 ;
        RECT 24.405 35.030 25.185 35.310 ;
        RECT 25.325 28.685 25.555 35.340 ;
        RECT 12.425 28.515 25.555 28.685 ;
        RECT 12.425 28.340 12.655 28.515 ;
        RECT 13.715 28.180 13.945 28.515 ;
        RECT 15.005 28.340 15.235 28.515 ;
        RECT 16.295 28.340 16.525 28.515 ;
        RECT 17.585 28.340 17.815 28.515 ;
        RECT 18.875 28.180 19.105 28.515 ;
        RECT 20.165 28.340 20.395 28.515 ;
        RECT 21.455 28.340 21.685 28.515 ;
        RECT 22.745 28.340 22.975 28.515 ;
        RECT 24.035 28.180 24.265 28.515 ;
        RECT 25.325 28.340 25.555 28.515 ;
        RECT 12.705 27.950 25.275 28.180 ;
        RECT 13.665 27.765 13.995 27.950 ;
        RECT 18.825 27.765 19.155 27.950 ;
        RECT 23.985 27.765 24.315 27.950 ;
        RECT 13.540 27.695 14.120 27.765 ;
        RECT 18.700 27.695 19.280 27.765 ;
        RECT 23.860 27.695 24.440 27.765 ;
        RECT 12.470 27.415 15.190 27.695 ;
        RECT 17.630 27.415 20.350 27.695 ;
        RECT 22.790 27.415 25.510 27.695 ;
        RECT 13.540 27.345 14.120 27.415 ;
        RECT 18.700 27.345 19.280 27.415 ;
        RECT 23.860 27.345 24.440 27.415 ;
        RECT 26.220 27.105 26.500 44.210 ;
        RECT 27.785 36.650 28.080 53.420 ;
        RECT 31.270 53.315 31.930 55.655 ;
        RECT 32.905 55.635 33.135 56.230 ;
        RECT 33.595 55.635 33.825 56.230 ;
        RECT 32.905 55.230 33.825 55.635 ;
        RECT 33.135 54.995 33.825 55.230 ;
        RECT 33.185 54.795 33.825 54.995 ;
        RECT 33.595 54.655 33.825 54.795 ;
        RECT 33.280 54.375 34.140 54.655 ;
        RECT 34.285 54.235 34.515 56.230 ;
        RECT 34.975 54.655 35.205 56.230 ;
        RECT 34.660 54.375 35.520 54.655 ;
        RECT 35.665 54.235 35.895 56.230 ;
        RECT 36.355 54.655 36.585 56.230 ;
        RECT 36.040 54.375 36.900 54.655 ;
        RECT 37.045 54.235 37.275 56.230 ;
        RECT 37.735 54.655 37.965 56.230 ;
        RECT 37.420 54.375 38.280 54.655 ;
        RECT 38.425 54.235 38.655 56.230 ;
        RECT 39.115 54.655 39.345 56.230 ;
        RECT 39.805 55.995 40.035 56.230 ;
        RECT 40.495 55.995 40.725 56.435 ;
        RECT 41.185 55.995 41.415 56.230 ;
        RECT 39.805 55.825 41.415 55.995 ;
        RECT 41.660 55.905 42.385 57.085 ;
        RECT 39.805 55.025 40.035 55.825 ;
        RECT 40.495 55.025 40.725 55.825 ;
        RECT 41.185 55.230 41.415 55.825 ;
        RECT 39.805 54.795 41.135 55.025 ;
        RECT 38.800 54.375 39.660 54.655 ;
        RECT 39.805 54.235 40.035 54.795 ;
        RECT 33.970 53.955 34.830 54.235 ;
        RECT 35.350 53.955 36.210 54.235 ;
        RECT 36.730 53.955 37.590 54.235 ;
        RECT 38.110 53.955 38.970 54.235 ;
        RECT 39.490 53.955 40.350 54.235 ;
        RECT 42.860 53.315 43.460 62.085 ;
        RECT 31.270 52.705 43.460 53.315 ;
        RECT 26.640 35.870 28.080 36.650 ;
        RECT 11.480 26.795 26.500 27.105 ;
        RECT 18.905 26.555 19.075 26.795 ;
        RECT 17.530 26.260 19.075 26.555 ;
        RECT 28.480 26.375 51.100 26.655 ;
        RECT 12.385 23.130 12.575 23.330 ;
        RECT 12.125 22.850 12.835 23.130 ;
        RECT 12.385 21.870 12.575 22.850 ;
        RECT 12.745 22.010 13.505 22.290 ;
        RECT 10.835 21.640 11.545 21.870 ;
        RECT 12.125 21.640 12.835 21.870 ;
        RECT 7.660 16.700 10.185 19.955 ;
        RECT 10.430 18.065 10.660 21.480 ;
        RECT 11.095 18.065 11.285 21.640 ;
        RECT 11.720 18.065 11.950 21.480 ;
        RECT 10.430 17.895 11.950 18.065 ;
        RECT 7.660 12.940 9.310 16.700 ;
        RECT 10.430 14.480 10.660 17.895 ;
        RECT 11.095 14.320 11.285 17.895 ;
        RECT 10.835 14.090 11.545 14.320 ;
        RECT 11.720 13.385 11.950 17.895 ;
        RECT 13.010 18.065 13.240 22.010 ;
        RECT 13.415 21.640 14.125 21.870 ;
        RECT 16.645 21.640 17.355 21.870 ;
        RECT 13.675 18.065 13.865 21.640 ;
        RECT 14.300 18.065 14.530 21.480 ;
        RECT 13.010 17.895 14.530 18.065 ;
        RECT 13.010 14.480 13.240 17.895 ;
        RECT 13.675 14.320 13.865 17.895 ;
        RECT 14.300 14.480 14.530 17.895 ;
        RECT 16.240 18.065 16.470 21.480 ;
        RECT 16.905 18.065 17.095 21.640 ;
        RECT 17.530 18.065 17.760 26.260 ;
        RECT 18.820 23.890 28.060 24.100 ;
        RECT 18.195 23.130 18.385 23.330 ;
        RECT 17.935 22.850 18.645 23.130 ;
        RECT 18.195 21.870 18.385 22.850 ;
        RECT 17.935 21.640 18.645 21.870 ;
        RECT 16.240 17.895 17.760 18.065 ;
        RECT 16.240 14.480 16.470 17.895 ;
        RECT 16.905 14.320 17.095 17.895 ;
        RECT 17.530 14.480 17.760 17.895 ;
        RECT 18.820 18.065 19.050 23.890 ;
        RECT 23.075 23.470 23.835 23.750 ;
        RECT 19.225 21.640 19.935 21.870 ;
        RECT 22.455 21.640 23.165 21.870 ;
        RECT 19.485 18.065 19.675 21.640 ;
        RECT 20.110 18.065 20.340 21.480 ;
        RECT 18.820 17.895 20.340 18.065 ;
        RECT 18.820 14.480 19.050 17.895 ;
        RECT 19.485 14.320 19.675 17.895 ;
        RECT 20.110 14.480 20.340 17.895 ;
        RECT 22.050 18.065 22.280 21.480 ;
        RECT 22.715 18.065 22.905 21.640 ;
        RECT 23.340 18.065 23.570 23.470 ;
        RECT 24.005 23.130 24.195 23.330 ;
        RECT 23.745 22.850 24.455 23.130 ;
        RECT 24.005 21.870 24.195 22.850 ;
        RECT 27.830 21.895 28.060 23.890 ;
        RECT 23.745 21.640 24.455 21.870 ;
        RECT 25.035 21.640 25.745 21.870 ;
        RECT 22.050 17.895 23.570 18.065 ;
        RECT 22.050 14.480 22.280 17.895 ;
        RECT 22.715 14.320 22.905 17.895 ;
        RECT 23.340 14.480 23.570 17.895 ;
        RECT 24.630 18.065 24.860 21.480 ;
        RECT 25.295 18.065 25.485 21.640 ;
        RECT 27.565 21.615 28.325 21.895 ;
        RECT 25.920 18.065 26.150 21.480 ;
        RECT 27.565 21.195 28.325 21.475 ;
        RECT 24.630 17.895 26.150 18.065 ;
        RECT 12.125 14.090 12.835 14.320 ;
        RECT 13.415 14.090 14.125 14.320 ;
        RECT 16.645 14.090 17.355 14.320 ;
        RECT 17.935 14.090 18.645 14.320 ;
        RECT 19.225 14.090 19.935 14.320 ;
        RECT 22.455 14.090 23.165 14.320 ;
        RECT 23.745 14.090 24.455 14.320 ;
        RECT 16.890 13.485 20.145 13.905 ;
        RECT 21.350 13.485 24.050 13.905 ;
        RECT 24.630 13.900 24.860 17.895 ;
        RECT 25.295 14.320 25.485 17.895 ;
        RECT 25.920 14.480 26.150 17.895 ;
        RECT 27.830 16.715 28.060 21.195 ;
        RECT 27.565 16.435 28.325 16.715 ;
        RECT 25.035 14.090 25.745 14.320 ;
        RECT 28.480 13.900 28.700 26.375 ;
        RECT 29.300 25.955 30.060 26.235 ;
        RECT 31.880 25.955 32.640 26.235 ;
        RECT 29.565 24.190 29.795 25.955 ;
        RECT 29.970 25.585 30.680 25.815 ;
        RECT 31.260 25.585 31.970 25.815 ;
        RECT 30.230 24.190 30.420 25.585 ;
        RECT 30.855 24.190 31.085 25.425 ;
        RECT 31.520 24.190 31.710 25.585 ;
        RECT 32.145 24.190 32.375 25.955 ;
        RECT 32.550 25.585 33.260 25.815 ;
        RECT 29.565 24.020 32.375 24.190 ;
        RECT 29.565 22.425 29.795 24.020 ;
        RECT 30.230 22.265 30.420 24.020 ;
        RECT 30.855 22.425 31.085 24.020 ;
        RECT 31.520 22.265 31.710 24.020 ;
        RECT 32.145 22.425 32.375 24.020 ;
        RECT 33.435 22.425 33.665 26.375 ;
        RECT 34.460 25.955 35.220 26.235 ;
        RECT 33.840 25.585 34.550 25.815 ;
        RECT 34.725 22.425 34.955 25.955 ;
        RECT 35.130 25.585 35.840 25.815 ;
        RECT 36.015 22.425 36.245 26.375 ;
        RECT 37.040 25.955 37.800 26.235 ;
        RECT 36.420 25.585 37.130 25.815 ;
        RECT 37.305 22.425 37.535 25.955 ;
        RECT 37.710 25.585 38.420 25.815 ;
        RECT 38.595 22.425 38.825 26.375 ;
        RECT 39.620 25.955 40.380 26.235 ;
        RECT 39.000 25.585 39.710 25.815 ;
        RECT 39.885 22.425 40.115 25.955 ;
        RECT 40.290 25.585 41.000 25.815 ;
        RECT 41.175 22.425 41.405 26.375 ;
        RECT 42.200 25.955 42.960 26.235 ;
        RECT 41.580 25.585 42.290 25.815 ;
        RECT 42.465 22.425 42.695 25.955 ;
        RECT 42.870 25.585 43.580 25.815 ;
        RECT 43.755 22.425 43.985 26.375 ;
        RECT 44.780 25.955 45.540 26.235 ;
        RECT 44.160 25.585 44.870 25.815 ;
        RECT 45.045 22.425 45.275 25.955 ;
        RECT 45.450 25.585 46.160 25.815 ;
        RECT 46.335 22.425 46.565 26.375 ;
        RECT 47.360 25.955 48.120 26.235 ;
        RECT 49.940 25.955 50.700 26.235 ;
        RECT 46.740 25.585 47.450 25.815 ;
        RECT 47.625 24.190 47.855 25.955 ;
        RECT 48.030 25.585 48.740 25.815 ;
        RECT 49.320 25.585 50.030 25.815 ;
        RECT 48.290 24.190 48.480 25.585 ;
        RECT 48.915 24.190 49.145 25.425 ;
        RECT 49.580 24.190 49.770 25.585 ;
        RECT 50.205 24.190 50.435 25.955 ;
        RECT 47.625 24.020 50.435 24.190 ;
        RECT 47.625 22.425 47.855 24.020 ;
        RECT 48.290 22.265 48.480 24.020 ;
        RECT 48.915 22.425 49.145 24.020 ;
        RECT 49.580 22.265 49.770 24.020 ;
        RECT 50.205 22.425 50.435 24.020 ;
        RECT 29.970 22.035 30.680 22.265 ;
        RECT 31.260 22.035 31.970 22.265 ;
        RECT 32.550 22.035 33.260 22.265 ;
        RECT 33.840 22.035 34.550 22.265 ;
        RECT 35.130 22.035 35.840 22.265 ;
        RECT 36.420 22.035 37.130 22.265 ;
        RECT 37.710 22.035 38.420 22.265 ;
        RECT 39.000 22.035 39.710 22.265 ;
        RECT 40.290 22.035 41.000 22.265 ;
        RECT 41.580 22.035 42.290 22.265 ;
        RECT 42.870 22.035 43.580 22.265 ;
        RECT 44.160 22.035 44.870 22.265 ;
        RECT 45.450 22.035 46.160 22.265 ;
        RECT 46.740 22.035 47.450 22.265 ;
        RECT 48.030 22.035 48.740 22.265 ;
        RECT 49.320 22.035 50.030 22.265 ;
        RECT 31.880 21.615 32.640 21.895 ;
        RECT 31.260 21.195 31.970 21.475 ;
        RECT 28.970 18.230 29.250 21.140 ;
        RECT 31.520 21.055 31.710 21.195 ;
        RECT 29.970 20.825 30.680 21.055 ;
        RECT 31.260 20.825 31.970 21.055 ;
        RECT 29.565 19.430 29.795 20.665 ;
        RECT 30.230 19.430 30.420 20.825 ;
        RECT 30.855 19.430 31.085 20.665 ;
        RECT 29.565 19.260 31.085 19.430 ;
        RECT 28.900 17.135 29.380 18.230 ;
        RECT 29.565 17.665 29.795 19.260 ;
        RECT 30.230 17.505 30.420 19.260 ;
        RECT 29.970 17.275 30.680 17.505 ;
        RECT 30.855 17.135 31.085 19.260 ;
        RECT 32.145 17.665 32.375 21.615 ;
        RECT 32.810 21.475 33.000 22.035 ;
        RECT 34.100 21.475 34.290 22.035 ;
        RECT 34.460 21.615 35.220 21.895 ;
        RECT 32.550 21.195 33.260 21.475 ;
        RECT 33.840 21.195 34.550 21.475 ;
        RECT 32.810 21.055 33.000 21.195 ;
        RECT 34.100 21.055 34.290 21.195 ;
        RECT 32.550 20.825 33.260 21.055 ;
        RECT 33.840 20.825 34.550 21.055 ;
        RECT 31.260 17.275 31.970 17.505 ;
        RECT 32.550 17.275 33.260 17.505 ;
        RECT 33.435 17.135 33.665 20.665 ;
        RECT 34.725 17.665 34.955 21.615 ;
        RECT 35.390 21.475 35.580 22.035 ;
        RECT 36.680 21.475 36.870 22.035 ;
        RECT 37.040 21.615 37.800 21.895 ;
        RECT 35.130 21.195 35.840 21.475 ;
        RECT 36.420 21.195 37.130 21.475 ;
        RECT 35.390 21.055 35.580 21.195 ;
        RECT 36.680 21.055 36.870 21.195 ;
        RECT 35.130 20.825 35.840 21.055 ;
        RECT 36.420 20.825 37.130 21.055 ;
        RECT 33.840 17.275 34.550 17.505 ;
        RECT 35.130 17.275 35.840 17.505 ;
        RECT 36.015 17.135 36.245 20.665 ;
        RECT 37.305 17.665 37.535 21.615 ;
        RECT 37.970 21.475 38.160 22.035 ;
        RECT 39.260 21.475 39.450 22.035 ;
        RECT 40.550 21.475 40.740 22.035 ;
        RECT 41.840 21.475 42.030 22.035 ;
        RECT 42.200 21.615 42.960 21.895 ;
        RECT 37.710 21.195 38.420 21.475 ;
        RECT 39.000 21.195 39.710 21.475 ;
        RECT 40.290 21.195 41.000 21.475 ;
        RECT 41.580 21.195 42.290 21.475 ;
        RECT 37.970 21.055 38.160 21.195 ;
        RECT 39.260 21.055 39.450 21.195 ;
        RECT 40.550 21.055 40.740 21.195 ;
        RECT 41.840 21.055 42.030 21.195 ;
        RECT 37.710 20.825 38.420 21.055 ;
        RECT 39.000 20.825 41.000 21.055 ;
        RECT 41.580 20.825 42.290 21.055 ;
        RECT 36.420 17.275 37.130 17.505 ;
        RECT 37.710 17.275 38.420 17.505 ;
        RECT 38.595 17.135 38.825 20.665 ;
        RECT 39.885 17.505 40.115 20.825 ;
        RECT 39.000 17.275 41.000 17.505 ;
        RECT 41.175 17.135 41.405 20.665 ;
        RECT 42.465 17.665 42.695 21.615 ;
        RECT 43.130 21.475 43.320 22.035 ;
        RECT 44.420 21.475 44.610 22.035 ;
        RECT 44.780 21.615 45.540 21.895 ;
        RECT 42.870 21.195 43.580 21.475 ;
        RECT 44.160 21.195 44.870 21.475 ;
        RECT 43.130 21.055 43.320 21.195 ;
        RECT 44.420 21.055 44.610 21.195 ;
        RECT 42.870 20.825 43.580 21.055 ;
        RECT 44.160 20.825 44.870 21.055 ;
        RECT 41.580 17.275 42.290 17.505 ;
        RECT 42.870 17.275 43.580 17.505 ;
        RECT 43.755 17.135 43.985 20.665 ;
        RECT 45.045 17.665 45.275 21.615 ;
        RECT 45.710 21.475 45.900 22.035 ;
        RECT 47.000 21.475 47.190 22.035 ;
        RECT 47.360 21.615 48.120 21.895 ;
        RECT 45.450 21.195 46.160 21.475 ;
        RECT 46.740 21.195 47.450 21.475 ;
        RECT 45.710 21.055 45.900 21.195 ;
        RECT 47.000 21.055 47.190 21.195 ;
        RECT 45.450 20.825 46.160 21.055 ;
        RECT 46.740 20.825 47.450 21.055 ;
        RECT 44.160 17.275 44.870 17.505 ;
        RECT 45.450 17.275 46.160 17.505 ;
        RECT 46.335 17.135 46.565 20.665 ;
        RECT 47.625 17.665 47.855 21.615 ;
        RECT 48.030 21.195 48.740 21.475 ;
        RECT 48.290 21.055 48.480 21.195 ;
        RECT 48.030 20.825 48.740 21.055 ;
        RECT 49.320 20.825 50.030 21.055 ;
        RECT 48.915 19.430 49.145 20.665 ;
        RECT 49.580 19.430 49.770 20.825 ;
        RECT 50.205 19.430 50.435 20.665 ;
        RECT 48.915 19.260 50.435 19.430 ;
        RECT 46.740 17.275 47.450 17.505 ;
        RECT 48.030 17.275 48.740 17.505 ;
        RECT 48.915 17.135 49.145 19.260 ;
        RECT 49.580 17.505 49.770 19.260 ;
        RECT 50.205 17.665 50.435 19.260 ;
        RECT 50.750 18.230 51.030 21.140 ;
        RECT 49.320 17.275 50.030 17.505 ;
        RECT 50.620 17.135 51.100 18.230 ;
        RECT 28.845 16.855 30.325 17.135 ;
        RECT 30.590 16.855 31.350 17.135 ;
        RECT 31.880 16.855 32.640 17.135 ;
        RECT 33.170 16.855 33.930 17.135 ;
        RECT 34.460 16.855 35.220 17.135 ;
        RECT 35.750 16.855 36.510 17.135 ;
        RECT 37.040 16.855 37.800 17.135 ;
        RECT 38.330 16.855 39.090 17.135 ;
        RECT 39.620 16.855 40.380 17.135 ;
        RECT 40.910 16.855 41.670 17.135 ;
        RECT 42.200 16.855 42.960 17.135 ;
        RECT 43.490 16.855 44.250 17.135 ;
        RECT 44.780 16.855 45.540 17.135 ;
        RECT 46.070 16.855 46.830 17.135 ;
        RECT 47.360 16.855 48.120 17.135 ;
        RECT 48.650 16.855 49.410 17.135 ;
        RECT 49.675 16.855 51.155 17.135 ;
        RECT 28.900 16.800 29.380 16.855 ;
        RECT 29.970 16.065 30.680 16.295 ;
        RECT 24.630 13.620 28.700 13.900 ;
        RECT 11.455 13.105 12.215 13.385 ;
        RECT 17.285 12.940 17.510 13.485 ;
        RECT 22.650 12.940 22.875 13.485 ;
        RECT 26.620 12.940 27.400 13.475 ;
        RECT 7.660 12.555 27.400 12.940 ;
        RECT 28.480 12.375 28.700 13.620 ;
        RECT 29.565 14.670 29.795 15.905 ;
        RECT 30.230 14.670 30.420 16.065 ;
        RECT 30.855 14.670 31.085 16.855 ;
        RECT 31.260 16.065 31.970 16.295 ;
        RECT 31.520 14.670 31.710 16.065 ;
        RECT 32.145 14.670 32.375 16.855 ;
        RECT 32.550 16.435 33.260 16.715 ;
        RECT 33.840 16.435 34.550 16.715 ;
        RECT 32.810 16.295 33.000 16.435 ;
        RECT 34.100 16.295 34.290 16.435 ;
        RECT 32.550 16.065 33.260 16.295 ;
        RECT 33.840 16.065 34.550 16.295 ;
        RECT 29.565 14.500 32.375 14.670 ;
        RECT 29.565 12.905 29.795 14.500 ;
        RECT 30.230 12.745 30.420 14.500 ;
        RECT 30.855 12.905 31.085 14.500 ;
        RECT 31.520 12.745 31.710 14.500 ;
        RECT 32.145 12.905 32.375 14.500 ;
        RECT 29.970 12.515 30.680 12.745 ;
        RECT 31.260 12.515 31.970 12.745 ;
        RECT 32.550 12.515 33.260 12.745 ;
        RECT 33.435 12.375 33.665 15.905 ;
        RECT 34.725 12.905 34.955 16.855 ;
        RECT 35.130 16.435 35.840 16.715 ;
        RECT 36.420 16.435 37.130 16.715 ;
        RECT 35.390 16.295 35.580 16.435 ;
        RECT 36.680 16.295 36.870 16.435 ;
        RECT 35.130 16.065 35.840 16.295 ;
        RECT 36.420 16.065 37.130 16.295 ;
        RECT 33.840 12.515 34.550 12.745 ;
        RECT 35.130 12.515 35.840 12.745 ;
        RECT 36.015 12.375 36.245 15.905 ;
        RECT 37.305 12.905 37.535 16.855 ;
        RECT 37.710 16.435 38.420 16.715 ;
        RECT 39.000 16.435 39.710 16.715 ;
        RECT 37.970 16.295 38.160 16.435 ;
        RECT 39.260 16.295 39.450 16.435 ;
        RECT 37.710 16.065 38.420 16.295 ;
        RECT 39.000 16.065 39.710 16.295 ;
        RECT 36.420 12.515 37.130 12.745 ;
        RECT 37.710 12.515 38.420 12.745 ;
        RECT 38.595 12.375 38.825 15.905 ;
        RECT 39.885 12.905 40.115 16.855 ;
        RECT 40.290 16.435 41.000 16.715 ;
        RECT 41.580 16.435 42.290 16.715 ;
        RECT 40.550 16.295 40.740 16.435 ;
        RECT 41.840 16.295 42.030 16.435 ;
        RECT 40.290 16.065 41.000 16.295 ;
        RECT 41.580 16.065 42.290 16.295 ;
        RECT 39.000 12.515 39.710 12.745 ;
        RECT 40.290 12.515 41.000 12.745 ;
        RECT 41.175 12.375 41.405 15.905 ;
        RECT 42.465 12.905 42.695 16.855 ;
        RECT 42.870 16.435 43.580 16.715 ;
        RECT 44.160 16.435 44.870 16.715 ;
        RECT 43.130 16.295 43.320 16.435 ;
        RECT 44.420 16.295 44.610 16.435 ;
        RECT 42.870 16.065 43.580 16.295 ;
        RECT 44.160 16.065 44.870 16.295 ;
        RECT 41.580 12.515 42.290 12.745 ;
        RECT 42.870 12.515 43.580 12.745 ;
        RECT 43.755 12.375 43.985 15.905 ;
        RECT 45.045 12.905 45.275 16.855 ;
        RECT 45.450 16.435 46.160 16.715 ;
        RECT 46.740 16.435 47.450 16.715 ;
        RECT 45.710 16.295 45.900 16.435 ;
        RECT 47.000 16.295 47.190 16.435 ;
        RECT 45.450 16.065 46.160 16.295 ;
        RECT 46.740 16.065 47.450 16.295 ;
        RECT 44.160 12.515 44.870 12.745 ;
        RECT 45.450 12.515 46.160 12.745 ;
        RECT 46.335 12.375 46.565 15.905 ;
        RECT 47.625 14.670 47.855 16.855 ;
        RECT 48.030 16.065 48.740 16.295 ;
        RECT 48.290 14.670 48.480 16.065 ;
        RECT 48.915 14.670 49.145 16.855 ;
        RECT 50.620 16.800 51.100 16.855 ;
        RECT 49.320 16.065 50.030 16.295 ;
        RECT 49.580 14.670 49.770 16.065 ;
        RECT 50.205 14.670 50.435 15.905 ;
        RECT 47.625 14.500 50.435 14.670 ;
        RECT 47.625 12.905 47.855 14.500 ;
        RECT 48.290 12.745 48.480 14.500 ;
        RECT 48.915 12.905 49.145 14.500 ;
        RECT 49.580 12.745 49.770 14.500 ;
        RECT 50.205 12.905 50.435 14.500 ;
        RECT 46.740 12.515 47.450 12.745 ;
        RECT 48.030 12.515 48.740 12.745 ;
        RECT 49.320 12.515 50.030 12.745 ;
        RECT 28.480 12.095 51.100 12.375 ;
      LAYER met2 ;
        RECT 1.000 65.650 31.280 66.890 ;
        RECT 53.510 65.940 54.250 66.900 ;
        RECT 29.100 64.515 94.750 64.795 ;
        RECT 8.530 61.355 26.220 61.595 ;
        RECT 8.530 60.635 9.310 61.355 ;
        RECT 13.055 61.005 14.550 61.355 ;
        RECT 18.215 61.005 19.710 61.355 ;
        RECT 23.375 61.005 24.870 61.355 ;
        RECT 26.640 54.090 26.920 62.180 ;
        RECT 10.640 53.810 26.920 54.090 ;
        RECT 7.230 31.000 8.830 31.960 ;
        RECT 9.475 27.345 9.755 52.830 ;
        RECT 10.640 35.310 10.920 53.810 ;
        RECT 27.060 53.670 27.340 62.185 ;
        RECT 12.180 53.390 27.340 53.670 ;
        RECT 12.705 52.970 26.920 53.250 ;
        RECT 11.060 52.550 25.800 52.830 ;
        RECT 11.060 35.730 11.340 52.550 ;
        RECT 26.640 36.150 26.920 52.970 ;
        RECT 12.180 35.870 26.920 36.150 ;
        RECT 11.060 35.450 25.275 35.730 ;
        RECT 10.640 35.030 25.800 35.310 ;
        RECT 27.060 34.890 27.340 53.390 ;
        RECT 12.180 34.610 27.340 34.890 ;
        RECT 27.480 60.095 27.760 62.175 ;
        RECT 29.100 60.095 29.740 64.515 ;
        RECT 27.480 59.845 29.740 60.095 ;
        RECT 27.480 54.235 27.760 59.845 ;
        RECT 29.100 54.745 29.740 59.845 ;
        RECT 28.140 54.235 29.740 54.745 ;
        RECT 30.500 64.095 42.290 64.375 ;
        RECT 30.500 63.775 31.280 64.095 ;
        RECT 93.910 63.835 94.750 64.515 ;
        RECT 30.500 61.945 31.125 63.775 ;
        RECT 30.500 61.665 42.280 61.945 ;
        RECT 30.500 57.085 31.125 61.665 ;
        RECT 30.500 56.805 42.310 57.085 ;
        RECT 30.500 54.655 31.125 56.805 ;
        RECT 30.500 54.375 42.205 54.655 ;
        RECT 27.480 53.955 42.330 54.235 ;
        RECT 27.480 53.925 29.100 53.955 ;
        RECT 13.055 27.345 14.550 27.695 ;
        RECT 18.215 27.345 19.710 27.695 ;
        RECT 23.375 27.345 24.870 27.695 ;
        RECT 8.530 27.105 26.500 27.345 ;
        RECT 8.530 26.385 9.310 27.105 ;
        RECT 9.475 24.105 9.755 27.105 ;
        RECT 27.480 26.655 27.760 53.925 ;
        RECT 28.140 53.830 29.100 53.925 ;
        RECT 29.935 53.420 114.070 53.700 ;
        RECT 113.230 52.740 114.070 53.420 ;
        RECT 6.900 23.675 9.755 24.105 ;
        RECT 23.340 26.375 27.760 26.655 ;
        RECT 23.340 23.750 23.570 26.375 ;
        RECT 27.050 25.955 51.760 26.235 ;
        RECT 6.900 10.285 7.140 23.675 ;
        RECT 23.075 23.470 23.835 23.750 ;
        RECT 25.530 23.330 26.370 23.555 ;
        RECT 10.210 22.595 26.370 23.330 ;
        RECT 7.280 22.010 13.505 22.290 ;
        RECT 7.280 10.670 7.520 22.010 ;
        RECT 27.050 17.135 27.400 25.955 ;
        RECT 27.565 21.615 51.100 21.895 ;
        RECT 27.565 21.195 51.100 21.475 ;
        RECT 27.050 16.855 52.825 17.135 ;
        RECT 27.050 13.475 27.400 16.855 ;
        RECT 27.565 16.435 51.100 16.715 ;
        RECT 11.455 13.105 26.110 13.385 ;
        RECT 25.840 12.335 26.110 13.105 ;
        RECT 26.620 12.555 27.400 13.475 ;
        RECT 27.830 12.335 28.060 16.435 ;
        RECT 25.840 12.100 28.060 12.335 ;
        RECT 7.280 10.425 153.145 10.670 ;
        RECT 6.900 10.040 133.825 10.285 ;
        RECT 132.985 1.570 133.825 10.040 ;
        RECT 152.305 1.570 153.145 10.425 ;
      LAYER met3 ;
        RECT 1.000 65.770 2.695 66.730 ;
        RECT 53.820 65.940 54.735 66.900 ;
        RECT 93.055 63.835 94.750 64.795 ;
        RECT 28.140 53.830 29.100 54.745 ;
        RECT 112.375 52.740 114.070 53.700 ;
        RECT 6.745 31.000 7.660 31.960 ;
        RECT 28.140 26.795 55.800 52.695 ;
        RECT 24.675 22.595 26.370 23.555 ;
        RECT 132.130 1.570 133.825 2.530 ;
        RECT 151.450 1.570 153.145 2.530 ;
      LAYER met4 ;
        RECT 28.140 53.830 29.100 54.745 ;
        RECT 54.250 54.210 55.080 66.900 ;
        RECT 93.055 63.835 94.750 64.795 ;
        RECT 6.000 31.000 7.230 31.960 ;
        RECT 28.160 26.855 28.640 53.830 ;
        RECT 44.880 53.225 55.080 54.210 ;
        RECT 44.880 52.300 50.550 53.225 ;
        RECT 30.295 27.190 55.405 52.300 ;
        RECT 24.675 23.110 26.370 23.555 ;
        RECT 24.675 22.810 27.770 23.110 ;
        RECT 24.675 22.595 26.370 22.810 ;
        RECT 27.470 11.665 27.770 22.810 ;
        RECT 93.850 11.665 94.750 63.835 ;
        RECT 112.375 52.740 114.070 53.700 ;
        RECT 113.170 11.665 114.070 52.740 ;
        RECT 138.310 11.665 138.610 224.760 ;
        RECT 27.470 11.365 138.610 11.665 ;
        RECT 93.850 1.000 94.750 11.365 ;
        RECT 113.170 1.000 114.070 11.365 ;
        RECT 132.130 1.570 133.825 2.530 ;
        RECT 151.450 1.570 153.145 2.530 ;
        RECT 132.490 1.000 133.390 1.570 ;
        RECT 151.810 1.000 152.710 1.570 ;
  END
END tt_um_lochidev_two_stage_opamp
END LIBRARY

