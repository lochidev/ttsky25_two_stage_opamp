* NGSPICE file created from ttsky25_two_stage_opamp.ext - technology: sky130A

.subckt ttsky25_two_stage_opamp VDD IBIAS VOUT VN VP EN VSS
X0 VSS.t126 VSS.t125 VSS.t126 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X1 VDD.t75 a_2479_7336.t18 VOUT.t25 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X2 VSS.t130 a_2080_2896.t5 a_2080_2896.t6 VSS.t33 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X3 VDD.t74 a_2479_7336.t19 VOUT.t18 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X4 VDD.t57 VDD.t56 VDD.t57 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X5 VSS.t138 a_2080_2896.t8 a_4920_2896.t23 VSS.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 VSS.t31 a_2080_2896.t9 a_4920_2896.t22 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X7 a_2479_7336.t15 a_2479_7336.t14 a_2479_7336.t15 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X8 VSS.t124 VSS.t123 VSS.t124 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X9 VDD.t55 VDD.t54 VDD.t55 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X10 VDD.t73 a_2479_7336.t20 VOUT.t21 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X11 VDD.t72 a_2479_7336.t21 VOUT.t24 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X12 a_4920_2896.t21 a_2080_2896.t10 VSS.t134 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X13 a_2479_7336.t13 a_2479_7336.t11 a_2479_7336.t12 VSS.t40 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X14 a_2479_7336.t6 VP.t0 a_2995_7336.t17 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X15 VSS.t38 a_2080_2896.t11 a_4920_2896.t20 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 VSS.t122 VSS.t121 VSS.t122 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X17 a_2995_7336.t9 VN.t0 a_2479_9004.t20 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X18 VDD.t71 a_2479_7336.t22 VOUT.t23 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X19 a_2479_9004.t19 VN.t1 a_2995_7336.t8 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X20 VSS.t120 VSS.t119 VSS.t120 VSS.t83 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X21 a_2479_9004.t12 a_2479_9004.t11 a_2479_9004.t12 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X22 VSS.t118 VSS.t117 VSS.t118 VSS.t52 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X23 a_4920_2896.t19 a_2080_2896.t12 VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X24 a_2479_9004.t10 a_2479_9004.t8 a_2479_9004.t9 VSS.t40 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X25 a_2479_9004.t18 VN.t2 a_2995_7336.t19 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X26 VSS.t50 a_2080_2896.t13 a_4920_2896.t18 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X27 VOUT.t16 a_2479_7336.t23 VDD.t70 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X28 VSS.t116 VSS.t115 VSS.t116 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X29 VDD.t53 VDD.t51 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X30 a_2995_7336.t16 VP.t1 a_2479_7336.t4 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X31 VSS.t114 VSS.t113 VSS.t114 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X32 a_3758_2896.t11 a_2080_2896.t14 VSS.t129 VSS.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X33 a_4920_2896.t17 a_2080_2896.t15 VSS.t55 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X34 a_2479_7336.t3 VP.t2 a_2995_7336.t15 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X35 a_3758_2896.t10 a_2080_2896.t16 VSS.t35 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X36 VOUT.t30 a_2479_7336.t24 VDD.t69 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X37 VSS.t137 a_2080_2896.t17 a_3758_2896.t9 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X38 a_4920_2896.t26 a_4920_2896.t25 a_4920_2896.t26 VSS.t24 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X39 a_4920_2896.t16 a_2080_2896.t18 VSS.t29 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X40 a_3758_2896.t8 a_2080_2896.t19 VSS.t133 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X41 a_3758_2896.t7 a_2080_2896.t20 VSS.t37 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X42 a_4920_2896.t24 EN.t0 VOUT.t0 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X43 a_2995_7336.t14 VP.t3 a_2479_7336.t5 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X44 VDD.t5 a_2479_9004.t6 a_2479_9004.t7 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X45 VOUT.t13 VOUT.t11 VOUT.t12 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X46 a_4920_2896.t15 a_2080_2896.t21 VSS.t44 VSS.t43 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X47 VDD.t50 VDD.t49 VDD.t50 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X48 VSS.t49 a_2080_2896.t22 a_4920_2896.t14 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X49 VDD.t48 VDD.t47 VDD.t48 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X50 VSS.t112 VSS.t111 VSS.t112 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X51 VDD.t68 a_2479_7336.t25 VOUT.t26 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X52 VSS.t110 VSS.t108 VSS.t109 VSS.t72 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X53 VSS.t107 VSS.t106 VSS.t107 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X54 VOUT.t10 VOUT.t8 VOUT.t9 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X55 VSS.t128 a_2080_2896.t23 a_4920_2896.t13 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X56 VOUT.t7 VOUT.t6 VOUT.t7 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X57 a_2995_7336.t1 VN.t3 a_2479_9004.t17 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X58 VDD.t67 a_2479_7336.t26 VOUT.t19 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X59 VSS.t105 VSS.t103 VSS.t104 VSS.t40 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X60 VDD.t46 VDD.t44 VDD.t45 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X61 a_2479_9004.t5 a_2479_9004.t4 VDD.t76 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X62 C1.t1 VOUT.t1 sky130_fd_pr__cap_mim_m3_1 l=25.5 w=25.5
X63 VDD.t66 a_2479_7336.t27 VOUT.t29 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X64 VSS.t54 a_2080_2896.t24 a_3758_2896.t6 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X65 a_4920_2896.t12 a_2080_2896.t25 VSS.t34 VSS.t33 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X66 VSS.t102 VSS.t101 VSS.t102 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X67 VOUT.t17 a_2479_7336.t28 VDD.t65 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X68 VDD.t10 a_2479_9004.t21 a_2479_7336.t10 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X69 VDD.t43 VDD.t42 VDD.t43 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X70 VSS.t100 VSS.t99 VSS.t100 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X71 VDD.t41 VDD.t40 VDD.t41 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X72 VOUT.t15 a_2479_7336.t29 VDD.t64 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X73 VSS.t136 a_2080_2896.t26 a_3758_2896.t5 VSS.t43 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X74 VSS.t98 VSS.t97 VSS.t98 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X75 VDD.t39 VDD.t38 VDD.t39 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X76 VSS.t96 VSS.t95 VSS.t96 VSS.t41 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X77 VDD.t37 VDD.t35 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X78 a_3758_2896.t4 a_2080_2896.t27 VSS.t28 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X79 VSS.t94 VSS.t93 VSS.t94 VSS.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X80 VSS.t92 VSS.t91 VSS.t92 VSS.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X81 VSS.t90 VSS.t89 VSS.t90 VSS.t83 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X82 a_2995_7336.t13 VP.t4 a_2479_7336.t1 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X83 VSS.t88 VSS.t87 VSS.t88 VSS.t52 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X84 a_4920_2896.t11 a_2080_2896.t28 VSS.t132 VSS.t45 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X85 a_2479_7336.t7 VP.t5 a_2995_7336.t12 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X86 a_2080_2896.t2 a_2080_2896.t0 a_2080_2896.t1 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X87 a_2479_7336.t8 a_2479_9004.t22 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X88 VSS.t131 a_2080_2896.t29 a_4920_2896.t10 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X89 a_2995_7336.t4 VN.t4 a_2479_9004.t16 VSS.t41 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X90 VOUT.t28 a_2479_7336.t30 VDD.t63 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X91 a_4920_2896.t9 a_2080_2896.t30 VSS.t42 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X92 a_2479_9004.t15 VN.t5 a_2995_7336.t0 VSS.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X93 VDD.t1 a_2479_9004.t23 a_2479_7336.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X94 VDD.t34 VDD.t32 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X95 VSS.t48 a_2080_2896.t31 a_4920_2896.t8 VSS.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X96 VOUT.t22 a_2479_7336.t31 VDD.t62 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X97 VSS.t127 a_2080_2896.t32 a_4920_2896.t7 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X98 a_2995_7336.t3 VN.t6 a_2479_9004.t14 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X99 VDD.t31 VDD.t29 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X100 a_4920_2896.t6 a_2080_2896.t33 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X101 a_2479_9004.t13 VN.t7 a_2995_7336.t18 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X102 VSS.t14 a_2080_2896.t34 a_4920_2896.t5 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X103 VSS.t86 VSS.t85 VSS.t86 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X104 a_2995_7336.t11 VP.t6 a_2479_7336.t16 VSS.t41 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X105 a_2479_7336.t17 VP.t7 a_2995_7336.t10 VSS.t17 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X106 VSS.t84 VSS.t82 VSS.t84 VSS.t83 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X107 VSS.t53 a_2080_2896.t35 a_3758_2896.t3 VSS.t52 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X108 VSS.t135 a_2080_2896.t36 a_3758_2896.t2 VSS.t45 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X109 VSS.t81 VSS.t79 VSS.t80 VSS.t72 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X110 a_3758_2896.t1 a_2080_2896.t37 VSS.t12 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X111 VDD.t6 a_2479_9004.t2 a_2479_9004.t3 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X112 VSS.t4 a_2080_2896.t38 a_3758_2896.t0 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X113 IBIAS.t1 IBIAS.t0 IBIAS.t1 VSS.t51 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X114 VSS.t78 VSS.t77 VSS.t78 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X115 VDD.t28 VDD.t27 VDD.t28 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X116 VSS.t10 a_2080_2896.t39 a_4920_2896.t4 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X117 VDD.t26 VDD.t24 VDD.t25 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X118 IBIAS.t2 EN.t1 a_2080_2896.t7 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X119 VSS.t76 VSS.t75 VSS.t76 VSS.t41 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X120 a_2479_7336.t2 a_2479_9004.t24 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X121 a_4920_2896.t3 a_2080_2896.t40 VSS.t58 VSS.t33 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X122 a_4920_2896.t2 a_2080_2896.t41 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X123 VOUT.t14 a_2479_7336.t32 VDD.t61 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X124 a_2479_7336.t9 C1.t0 VSS.t32 sky130_fd_pr__res_xhigh_po_1p41 l=14
X125 VDD.t23 VDD.t21 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X126 VDD.t20 VDD.t18 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X127 a_3758_2896.t14 a_3758_2896.t13 a_3758_2896.t14 VSS.t57 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X128 VOUT.t31 a_2479_7336.t33 VDD.t60 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X129 VOUT.t5 VOUT.t4 VOUT.t5 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X130 a_4920_2896.t1 a_2080_2896.t42 VSS.t56 VSS.t43 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X131 a_3758_2896.t12 EN.t2 a_2995_7336.t2 VSS.t21 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X132 VSS.t27 a_2080_2896.t43 a_4920_2896.t0 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X133 VOUT.t3 VOUT.t2 VOUT.t3 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X134 VOUT.t27 a_2479_7336.t34 VDD.t59 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X135 VSS.t74 VSS.t71 VSS.t73 VSS.t72 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X136 a_2995_7336.t7 a_2995_7336.t5 a_2995_7336.t6 VSS.t59 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X137 VDD.t17 VDD.t15 VDD.t17 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X138 VSS.t70 VSS.t69 VSS.t70 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X139 VDD.t14 VDD.t11 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X140 a_2080_2896.t4 a_2080_2896.t3 VSS.t39 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X141 VSS.t68 VSS.t66 VSS.t67 VSS.t40 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X142 VSS.t65 VSS.t64 VSS.t65 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X143 VDD.t58 a_2479_7336.t35 VOUT.t20 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X144 VSS.t63 VSS.t62 VSS.t63 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X145 a_2479_9004.t1 a_2479_9004.t0 VDD.t7 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X146 VSS.t61 VSS.t60 VSS.t61 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
R0 VSS.n2193 VSS.n2192 2542.66
R1 VSS.n561 VSS.n546 1321.06
R2 VSS.n559 VSS.n548 1321.06
R3 VSS.n2194 VSS.n525 1321.06
R4 VSS.n642 VSS.n531 1321.06
R5 VSS.n2012 VSS.n874 1268.91
R6 VSS.n2081 VSS.n900 1268.91
R7 VSS.n2016 VSS.n2015 1268.91
R8 VSS.n2037 VSS.n2036 1268.91
R9 VSS.n1722 VSS.n1658 1268.91
R10 VSS.n1808 VSS.n1410 1268.91
R11 VSS.n1681 VSS.n1655 1268.91
R12 VSS.n1765 VSS.n1422 1268.91
R13 VSS.n744 VSS.n702 1268.91
R14 VSS.n2127 VSS.n777 1268.91
R15 VSS.n857 VSS.n774 1268.91
R16 VSS.n2161 VSS.n696 1268.91
R17 VSS.n432 VSS.n219 1182
R18 VSS.n2554 VSS.n101 1182
R19 VSS.n430 VSS.n221 1182
R20 VSS.n2490 VSS.n106 1182
R21 VSS.n2190 VSS.n655 1182
R22 VSS.n1171 VSS.n940 1182
R23 VSS.n1726 VSS.n1433 1182
R24 VSS.n2096 VSS.n887 1182
R25 VSS.n1130 VSS.n954 996.588
R26 VSS.n2193 VSS.n524 614.067
R27 VSS.n1082 VSS.n966 602.588
R28 VSS.n1034 VSS.n978 602.588
R29 VSS.n608 VSS.n607 585
R30 VSS.n607 VSS.n480 585
R31 VSS.n606 VSS.n479 585
R32 VSS.n2255 VSS.n479 585
R33 VSS.n605 VSS.n604 585
R34 VSS.n604 VSS.n475 585
R35 VSS.n603 VSS.n474 585
R36 VSS.n2261 VSS.n474 585
R37 VSS.n602 VSS.n473 585
R38 VSS.n2262 VSS.n473 585
R39 VSS.n601 VSS.n472 585
R40 VSS.n2263 VSS.n472 585
R41 VSS.n600 VSS.n599 585
R42 VSS.n599 VSS.n468 585
R43 VSS.n598 VSS.n467 585
R44 VSS.n2269 VSS.n467 585
R45 VSS.n597 VSS.n466 585
R46 VSS.n2270 VSS.n466 585
R47 VSS.n596 VSS.n465 585
R48 VSS.n2271 VSS.n465 585
R49 VSS.n595 VSS.n594 585
R50 VSS.n594 VSS.n461 585
R51 VSS.n593 VSS.n460 585
R52 VSS.n2277 VSS.n460 585
R53 VSS.n592 VSS.n459 585
R54 VSS.n2278 VSS.n459 585
R55 VSS.n591 VSS.n458 585
R56 VSS.n2279 VSS.n458 585
R57 VSS.n590 VSS.n589 585
R58 VSS.n589 VSS.n454 585
R59 VSS.n588 VSS.n453 585
R60 VSS.n2285 VSS.n453 585
R61 VSS.n587 VSS.n452 585
R62 VSS.n2286 VSS.n452 585
R63 VSS.n586 VSS.n451 585
R64 VSS.n2287 VSS.n451 585
R65 VSS.n585 VSS.n584 585
R66 VSS.n584 VSS.n445 585
R67 VSS.n583 VSS.n444 585
R68 VSS.n2293 VSS.n444 585
R69 VSS.n582 VSS.n581 585
R70 VSS.n581 VSS.n443 585
R71 VSS.n580 VSS.n533 585
R72 VSS.n580 VSS.n579 585
R73 VSS.n570 VSS.n534 585
R74 VSS.n535 VSS.n534 585
R75 VSS.n572 VSS.n571 585
R76 VSS.n573 VSS.n572 585
R77 VSS.n569 VSS.n540 585
R78 VSS.n540 VSS.n539 585
R79 VSS.n568 VSS.n567 585
R80 VSS.n567 VSS.n566 585
R81 VSS.n542 VSS.n541 585
R82 VSS.n543 VSS.n542 585
R83 VSS.n559 VSS.n558 585
R84 VSS.n560 VSS.n559 585
R85 VSS.n557 VSS.n548 585
R86 VSS.n556 VSS.n555 585
R87 VSS.n553 VSS.n549 585
R88 VSS.n551 VSS.n550 585
R89 VSS.n546 VSS.n545 585
R90 VSS.n547 VSS.n546 585
R91 VSS.n562 VSS.n561 585
R92 VSS.n561 VSS.n560 585
R93 VSS.n563 VSS.n544 585
R94 VSS.n544 VSS.n543 585
R95 VSS.n565 VSS.n564 585
R96 VSS.n566 VSS.n565 585
R97 VSS.n538 VSS.n537 585
R98 VSS.n539 VSS.n538 585
R99 VSS.n575 VSS.n574 585
R100 VSS.n574 VSS.n573 585
R101 VSS.n576 VSS.n536 585
R102 VSS.n536 VSS.n535 585
R103 VSS.n578 VSS.n577 585
R104 VSS.n579 VSS.n578 585
R105 VSS.n448 VSS.n446 585
R106 VSS.n446 VSS.n443 585
R107 VSS.n2292 VSS.n2291 585
R108 VSS.n2293 VSS.n2292 585
R109 VSS.n2290 VSS.n447 585
R110 VSS.n447 VSS.n445 585
R111 VSS.n2289 VSS.n2288 585
R112 VSS.n2288 VSS.n2287 585
R113 VSS.n450 VSS.n449 585
R114 VSS.n2286 VSS.n450 585
R115 VSS.n2284 VSS.n2283 585
R116 VSS.n2285 VSS.n2284 585
R117 VSS.n2282 VSS.n455 585
R118 VSS.n455 VSS.n454 585
R119 VSS.n2281 VSS.n2280 585
R120 VSS.n2280 VSS.n2279 585
R121 VSS.n457 VSS.n456 585
R122 VSS.n2278 VSS.n457 585
R123 VSS.n2276 VSS.n2275 585
R124 VSS.n2277 VSS.n2276 585
R125 VSS.n2274 VSS.n462 585
R126 VSS.n462 VSS.n461 585
R127 VSS.n2273 VSS.n2272 585
R128 VSS.n2272 VSS.n2271 585
R129 VSS.n464 VSS.n463 585
R130 VSS.n2270 VSS.n464 585
R131 VSS.n2268 VSS.n2267 585
R132 VSS.n2269 VSS.n2268 585
R133 VSS.n2266 VSS.n469 585
R134 VSS.n469 VSS.n468 585
R135 VSS.n2265 VSS.n2264 585
R136 VSS.n2264 VSS.n2263 585
R137 VSS.n471 VSS.n470 585
R138 VSS.n2262 VSS.n471 585
R139 VSS.n2260 VSS.n2259 585
R140 VSS.n2261 VSS.n2260 585
R141 VSS.n2258 VSS.n476 585
R142 VSS.n476 VSS.n475 585
R143 VSS.n2257 VSS.n2256 585
R144 VSS.n2256 VSS.n2255 585
R145 VSS.n478 VSS.n477 585
R146 VSS.n480 VSS.n478 585
R147 VSS.n2194 VSS.n526 585
R148 VSS.n2197 VSS.n2196 585
R149 VSS.n529 VSS.n528 585
R150 VSS.n2193 VSS.n529 585
R151 VSS.n532 VSS.n530 585
R152 VSS.n642 VSS.n641 585
R153 VSS.n640 VSS.n531 585
R154 VSS.n531 VSS.n524 585
R155 VSS.n639 VSS.n523 585
R156 VSS.n2205 VSS.n523 585
R157 VSS.n638 VSS.n522 585
R158 VSS.n2206 VSS.n522 585
R159 VSS.n637 VSS.n521 585
R160 VSS.n2207 VSS.n521 585
R161 VSS.n636 VSS.n635 585
R162 VSS.n635 VSS.n517 585
R163 VSS.n634 VSS.n516 585
R164 VSS.n2213 VSS.n516 585
R165 VSS.n633 VSS.n515 585
R166 VSS.n2214 VSS.n515 585
R167 VSS.n632 VSS.n514 585
R168 VSS.n2215 VSS.n514 585
R169 VSS.n631 VSS.n630 585
R170 VSS.n630 VSS.n510 585
R171 VSS.n629 VSS.n509 585
R172 VSS.n2221 VSS.n509 585
R173 VSS.n628 VSS.n508 585
R174 VSS.n2222 VSS.n508 585
R175 VSS.n627 VSS.n507 585
R176 VSS.n2223 VSS.n507 585
R177 VSS.n626 VSS.n625 585
R178 VSS.n625 VSS.n503 585
R179 VSS.n624 VSS.n502 585
R180 VSS.n2229 VSS.n502 585
R181 VSS.n623 VSS.n501 585
R182 VSS.n2230 VSS.n501 585
R183 VSS.n622 VSS.n500 585
R184 VSS.n2231 VSS.n500 585
R185 VSS.n621 VSS.n620 585
R186 VSS.n620 VSS.n496 585
R187 VSS.n619 VSS.n495 585
R188 VSS.n2237 VSS.n495 585
R189 VSS.n618 VSS.n494 585
R190 VSS.n2238 VSS.n494 585
R191 VSS.n617 VSS.n493 585
R192 VSS.n2239 VSS.n493 585
R193 VSS.n616 VSS.n615 585
R194 VSS.n615 VSS.n489 585
R195 VSS.n614 VSS.n488 585
R196 VSS.n2245 VSS.n488 585
R197 VSS.n613 VSS.n487 585
R198 VSS.n2246 VSS.n487 585
R199 VSS.n612 VSS.n486 585
R200 VSS.n2247 VSS.n486 585
R201 VSS.n611 VSS.n610 585
R202 VSS.n610 VSS.n482 585
R203 VSS.n609 VSS.n481 585
R204 VSS.n2253 VSS.n481 585
R205 VSS.n2252 VSS.n2251 585
R206 VSS.n2253 VSS.n2252 585
R207 VSS.n2250 VSS.n483 585
R208 VSS.n483 VSS.n482 585
R209 VSS.n2249 VSS.n2248 585
R210 VSS.n2248 VSS.n2247 585
R211 VSS.n485 VSS.n484 585
R212 VSS.n2246 VSS.n485 585
R213 VSS.n2244 VSS.n2243 585
R214 VSS.n2245 VSS.n2244 585
R215 VSS.n2242 VSS.n490 585
R216 VSS.n490 VSS.n489 585
R217 VSS.n2241 VSS.n2240 585
R218 VSS.n2240 VSS.n2239 585
R219 VSS.n492 VSS.n491 585
R220 VSS.n2238 VSS.n492 585
R221 VSS.n2236 VSS.n2235 585
R222 VSS.n2237 VSS.n2236 585
R223 VSS.n2234 VSS.n497 585
R224 VSS.n497 VSS.n496 585
R225 VSS.n2233 VSS.n2232 585
R226 VSS.n2232 VSS.n2231 585
R227 VSS.n499 VSS.n498 585
R228 VSS.n2230 VSS.n499 585
R229 VSS.n2228 VSS.n2227 585
R230 VSS.n2229 VSS.n2228 585
R231 VSS.n2226 VSS.n504 585
R232 VSS.n504 VSS.n503 585
R233 VSS.n2225 VSS.n2224 585
R234 VSS.n2224 VSS.n2223 585
R235 VSS.n506 VSS.n505 585
R236 VSS.n2222 VSS.n506 585
R237 VSS.n2220 VSS.n2219 585
R238 VSS.n2221 VSS.n2220 585
R239 VSS.n2218 VSS.n511 585
R240 VSS.n511 VSS.n510 585
R241 VSS.n2217 VSS.n2216 585
R242 VSS.n2216 VSS.n2215 585
R243 VSS.n513 VSS.n512 585
R244 VSS.n2214 VSS.n513 585
R245 VSS.n2212 VSS.n2211 585
R246 VSS.n2213 VSS.n2212 585
R247 VSS.n2210 VSS.n518 585
R248 VSS.n518 VSS.n517 585
R249 VSS.n2209 VSS.n2208 585
R250 VSS.n2208 VSS.n2207 585
R251 VSS.n520 VSS.n519 585
R252 VSS.n2206 VSS.n520 585
R253 VSS.n2204 VSS.n2203 585
R254 VSS.n2205 VSS.n2204 585
R255 VSS.n2202 VSS.n525 585
R256 VSS.n525 VSS.n524 585
R257 VSS.n1171 VSS.n1170 585
R258 VSS.n1169 VSS.n951 585
R259 VSS.n1168 VSS.n950 585
R260 VSS.n1173 VSS.n950 585
R261 VSS.n1167 VSS.n1166 585
R262 VSS.n1165 VSS.n1164 585
R263 VSS.n1163 VSS.n1162 585
R264 VSS.n1161 VSS.n1160 585
R265 VSS.n1159 VSS.n1158 585
R266 VSS.n1157 VSS.n1156 585
R267 VSS.n1155 VSS.n1154 585
R268 VSS.n1153 VSS.n1152 585
R269 VSS.n1151 VSS.n1150 585
R270 VSS.n1149 VSS.n1148 585
R271 VSS.n1147 VSS.n1146 585
R272 VSS.n1145 VSS.n1144 585
R273 VSS.n1143 VSS.n1142 585
R274 VSS.n1141 VSS.n1140 585
R275 VSS.n1139 VSS.n1138 585
R276 VSS.n1137 VSS.n1136 585
R277 VSS.n1135 VSS.n949 585
R278 VSS.n1173 VSS.n949 585
R279 VSS.n1510 VSS.n1509 585
R280 VSS.n1508 VSS.n1507 585
R281 VSS.n1506 VSS.n1505 585
R282 VSS.n1504 VSS.n1503 585
R283 VSS.n1502 VSS.n1501 585
R284 VSS.n1500 VSS.n1499 585
R285 VSS.n1498 VSS.n1497 585
R286 VSS.n1496 VSS.n1495 585
R287 VSS.n1494 VSS.n1493 585
R288 VSS.n1492 VSS.n1491 585
R289 VSS.n1490 VSS.n1489 585
R290 VSS.n1488 VSS.n1487 585
R291 VSS.n1486 VSS.n1485 585
R292 VSS.n1484 VSS.n1483 585
R293 VSS.n1482 VSS.n1481 585
R294 VSS.n1480 VSS.n1479 585
R295 VSS.n1478 VSS.n1477 585
R296 VSS.n1476 VSS.n1475 585
R297 VSS.n1474 VSS.n1473 585
R298 VSS.n657 VSS.n655 585
R299 VSS.n2190 VSS.n2189 585
R300 VSS.n2191 VSS.n2190 585
R301 VSS.n658 VSS.n656 585
R302 VSS.n656 VSS.n654 585
R303 VSS.n2185 VSS.n2184 585
R304 VSS.n2184 VSS.n2183 585
R305 VSS.n661 VSS.n660 585
R306 VSS.n2182 VSS.n661 585
R307 VSS.n2180 VSS.n2179 585
R308 VSS.n2181 VSS.n2180 585
R309 VSS.n2178 VSS.n663 585
R310 VSS.n663 VSS.n662 585
R311 VSS.n1749 VSS.n665 585
R312 VSS.n1750 VSS.n1749 585
R313 VSS.n669 VSS.n667 585
R314 VSS.n671 VSS.n669 585
R315 VSS.n2174 VSS.n2173 585
R316 VSS.n2173 VSS.n2172 585
R317 VSS.n670 VSS.n668 585
R318 VSS.n2171 VSS.n670 585
R319 VSS.n1304 VSS.n1303 585
R320 VSS.n1303 VSS.n672 585
R321 VSS.n1306 VSS.n1305 585
R322 VSS.n1307 VSS.n1306 585
R323 VSS.n1309 VSS.n1302 585
R324 VSS.n1309 VSS.n1308 585
R325 VSS.n1311 VSS.n1310 585
R326 VSS.n1310 VSS.n681 585
R327 VSS.n1312 VSS.n1301 585
R328 VSS.n1301 VSS.n682 585
R329 VSS.n1314 VSS.n1313 585
R330 VSS.n1315 VSS.n1314 585
R331 VSS.n1317 VSS.n1299 585
R332 VSS.n1317 VSS.n1316 585
R333 VSS.n1908 VSS.n1907 585
R334 VSS.n1907 VSS.n1906 585
R335 VSS.n1318 VSS.n1300 585
R336 VSS.n1323 VSS.n1318 585
R337 VSS.n1321 VSS.n1320 585
R338 VSS.n1322 VSS.n1321 585
R339 VSS.n1192 VSS.n1191 585
R340 VSS.n1319 VSS.n1191 585
R341 VSS.n1920 VSS.n1919 585
R342 VSS.n1921 VSS.n1920 585
R343 VSS.n1193 VSS.n1190 585
R344 VSS.n1922 VSS.n1190 585
R345 VSS.n1926 VSS.n1925 585
R346 VSS.n1925 VSS.n1924 585
R347 VSS.n1927 VSS.n1188 585
R348 VSS.n1923 VSS.n1188 585
R349 VSS.n1929 VSS.n1928 585
R350 VSS.n1930 VSS.n1929 585
R351 VSS.n1186 VSS.n1185 585
R352 VSS.n1931 VSS.n1186 585
R353 VSS.n1934 VSS.n1933 585
R354 VSS.n1933 VSS.n1932 585
R355 VSS.n1935 VSS.n1184 585
R356 VSS.n1184 VSS.n859 585
R357 VSS.n1937 VSS.n1936 585
R358 VSS.n1937 VSS.n860 585
R359 VSS.n1938 VSS.n1182 585
R360 VSS.n1939 VSS.n1938 585
R361 VSS.n1942 VSS.n1941 585
R362 VSS.n1941 VSS.n1940 585
R363 VSS.n1183 VSS.n928 585
R364 VSS.n928 VSS.n926 585
R365 VSS.n1955 VSS.n1954 585
R366 VSS.n1956 VSS.n1955 585
R367 VSS.n1953 VSS.n929 585
R368 VSS.n929 VSS.n927 585
R369 VSS.n936 VSS.n931 585
R370 VSS.n937 VSS.n936 585
R371 VSS.n939 VSS.n935 585
R372 VSS.n939 VSS.n938 585
R373 VSS.n1177 VSS.n1176 585
R374 VSS.n1176 VSS.n1175 585
R375 VSS.n952 VSS.n940 585
R376 VSS.n1174 VSS.n940 585
R377 VSS.n1809 VSS.n1808 585
R378 VSS.n1806 VSS.n1411 585
R379 VSS.n1805 VSS.n1804 585
R380 VSS.n1805 VSS.n680 585
R381 VSS.n1803 VSS.n1412 585
R382 VSS.n1802 VSS.n1801 585
R383 VSS.n1799 VSS.n1413 585
R384 VSS.n1797 VSS.n1796 585
R385 VSS.n1795 VSS.n1414 585
R386 VSS.n1794 VSS.n1793 585
R387 VSS.n1791 VSS.n1415 585
R388 VSS.n1789 VSS.n1788 585
R389 VSS.n1787 VSS.n1416 585
R390 VSS.n1786 VSS.n1785 585
R391 VSS.n1783 VSS.n1417 585
R392 VSS.n1781 VSS.n1780 585
R393 VSS.n1779 VSS.n1418 585
R394 VSS.n1778 VSS.n1777 585
R395 VSS.n1775 VSS.n1419 585
R396 VSS.n1773 VSS.n1772 585
R397 VSS.n1771 VSS.n1420 585
R398 VSS.n1770 VSS.n1769 585
R399 VSS.n1767 VSS.n1421 585
R400 VSS.n1765 VSS.n1764 585
R401 VSS.n1423 VSS.n1422 585
R402 VSS.n1422 VSS.n673 585
R403 VSS.n1760 VSS.n1408 585
R404 VSS.n1813 VSS.n1408 585
R405 VSS.n1759 VSS.n1758 585
R406 VSS.n1758 VSS.n1406 585
R407 VSS.n1424 VSS.n1405 585
R408 VSS.n1825 VSS.n1405 585
R409 VSS.n1753 VSS.n1752 585
R410 VSS.n1752 VSS.n1751 585
R411 VSS.n1747 VSS.n1397 585
R412 VSS.n1831 VSS.n1397 585
R413 VSS.n1746 VSS.n1745 585
R414 VSS.n1745 VSS.n1744 585
R415 VSS.n1426 VSS.n1425 585
R416 VSS.n1742 VSS.n1426 585
R417 VSS.n1675 VSS.n1674 585
R418 VSS.n1674 VSS.n1432 585
R419 VSS.n1676 VSS.n1431 585
R420 VSS.n1736 VSS.n1431 585
R421 VSS.n1678 VSS.n1677 585
R422 VSS.n1677 VSS.n1657 585
R423 VSS.n1679 VSS.n1655 585
R424 VSS.n1723 VSS.n1655 585
R425 VSS.n1682 VSS.n1681 585
R426 VSS.n1683 VSS.n1673 585
R427 VSS.n1685 VSS.n1684 585
R428 VSS.n1687 VSS.n1671 585
R429 VSS.n1689 VSS.n1688 585
R430 VSS.n1690 VSS.n1670 585
R431 VSS.n1692 VSS.n1691 585
R432 VSS.n1694 VSS.n1668 585
R433 VSS.n1696 VSS.n1695 585
R434 VSS.n1697 VSS.n1667 585
R435 VSS.n1699 VSS.n1698 585
R436 VSS.n1701 VSS.n1665 585
R437 VSS.n1703 VSS.n1702 585
R438 VSS.n1704 VSS.n1664 585
R439 VSS.n1706 VSS.n1705 585
R440 VSS.n1708 VSS.n1662 585
R441 VSS.n1710 VSS.n1709 585
R442 VSS.n1711 VSS.n1661 585
R443 VSS.n1713 VSS.n1712 585
R444 VSS.n1715 VSS.n1660 585
R445 VSS.n1716 VSS.n1659 585
R446 VSS.n1719 VSS.n1718 585
R447 VSS.n1720 VSS.n1658 585
R448 VSS.n1658 VSS.n98 585
R449 VSS.n1722 VSS.n1721 585
R450 VSS.n1723 VSS.n1722 585
R451 VSS.n1430 VSS.n1429 585
R452 VSS.n1657 VSS.n1430 585
R453 VSS.n1738 VSS.n1737 585
R454 VSS.n1737 VSS.n1736 585
R455 VSS.n1739 VSS.n1428 585
R456 VSS.n1432 VSS.n1428 585
R457 VSS.n1741 VSS.n1740 585
R458 VSS.n1742 VSS.n1741 585
R459 VSS.n1401 VSS.n1399 585
R460 VSS.n1744 VSS.n1399 585
R461 VSS.n1830 VSS.n1829 585
R462 VSS.n1831 VSS.n1830 585
R463 VSS.n1828 VSS.n1400 585
R464 VSS.n1751 VSS.n1400 585
R465 VSS.n1827 VSS.n1826 585
R466 VSS.n1826 VSS.n1825 585
R467 VSS.n1403 VSS.n1402 585
R468 VSS.n1406 VSS.n1403 585
R469 VSS.n1812 VSS.n1811 585
R470 VSS.n1813 VSS.n1812 585
R471 VSS.n1810 VSS.n1410 585
R472 VSS.n1410 VSS.n673 585
R473 VSS.n2082 VSS.n2081 585
R474 VSS.n902 VSS.n901 585
R475 VSS.n2078 VSS.n2077 585
R476 VSS.n2079 VSS.n2078 585
R477 VSS.n2076 VSS.n913 585
R478 VSS.n2075 VSS.n2074 585
R479 VSS.n2073 VSS.n2072 585
R480 VSS.n2071 VSS.n2070 585
R481 VSS.n2069 VSS.n2068 585
R482 VSS.n918 VSS.n915 585
R483 VSS.n920 VSS.n919 585
R484 VSS.n2063 VSS.n2062 585
R485 VSS.n2061 VSS.n2060 585
R486 VSS.n2059 VSS.n2058 585
R487 VSS.n2057 VSS.n2056 585
R488 VSS.n2054 VSS.n2053 585
R489 VSS.n2052 VSS.n2051 585
R490 VSS.n2050 VSS.n2049 585
R491 VSS.n2048 VSS.n2047 585
R492 VSS.n2046 VSS.n2045 585
R493 VSS.n2044 VSS.n2043 585
R494 VSS.n2042 VSS.n2041 585
R495 VSS.n2040 VSS.n2039 585
R496 VSS.n2038 VSS.n2037 585
R497 VSS.n2036 VSS.n2035 585
R498 VSS.n2036 VSS.n899 585
R499 VSS.n2034 VSS.n898 585
R500 VSS.n2086 VSS.n898 585
R501 VSS.n2033 VSS.n897 585
R502 VSS.n2087 VSS.n897 585
R503 VSS.n2032 VSS.n896 585
R504 VSS.n2088 VSS.n896 585
R505 VSS.n2031 VSS.n2030 585
R506 VSS.n2030 VSS.n890 585
R507 VSS.n2029 VSS.n889 585
R508 VSS.n2094 VSS.n889 585
R509 VSS.n2028 VSS.n2027 585
R510 VSS.n2027 VSS.n888 585
R511 VSS.n2026 VSS.n2023 585
R512 VSS.n2026 VSS.n2025 585
R513 VSS.n2022 VSS.n880 585
R514 VSS.n2104 VSS.n880 585
R515 VSS.n2021 VSS.n2020 585
R516 VSS.n2020 VSS.n2019 585
R517 VSS.n2018 VSS.n872 585
R518 VSS.n2110 VSS.n872 585
R519 VSS.n2017 VSS.n2016 585
R520 VSS.n2016 VSS.n871 585
R521 VSS.n2015 VSS.n924 585
R522 VSS.n1971 VSS.n925 585
R523 VSS.n1973 VSS.n1972 585
R524 VSS.n1975 VSS.n1974 585
R525 VSS.n1977 VSS.n1976 585
R526 VSS.n1979 VSS.n1978 585
R527 VSS.n1981 VSS.n1980 585
R528 VSS.n1983 VSS.n1982 585
R529 VSS.n1985 VSS.n1984 585
R530 VSS.n1987 VSS.n1986 585
R531 VSS.n1989 VSS.n1988 585
R532 VSS.n1991 VSS.n1990 585
R533 VSS.n1993 VSS.n1992 585
R534 VSS.n1995 VSS.n1994 585
R535 VSS.n1997 VSS.n1996 585
R536 VSS.n1999 VSS.n1998 585
R537 VSS.n2001 VSS.n2000 585
R538 VSS.n2003 VSS.n2002 585
R539 VSS.n2005 VSS.n2004 585
R540 VSS.n2007 VSS.n2006 585
R541 VSS.n2009 VSS.n2008 585
R542 VSS.n2010 VSS.n1970 585
R543 VSS.n2012 VSS.n2011 585
R544 VSS.n2013 VSS.n2012 585
R545 VSS.n876 VSS.n874 585
R546 VSS.n874 VSS.n871 585
R547 VSS.n2109 VSS.n2108 585
R548 VSS.n2110 VSS.n2109 585
R549 VSS.n2107 VSS.n875 585
R550 VSS.n2019 VSS.n875 585
R551 VSS.n2106 VSS.n2105 585
R552 VSS.n2105 VSS.n2104 585
R553 VSS.n878 VSS.n877 585
R554 VSS.n2025 VSS.n878 585
R555 VSS.n893 VSS.n891 585
R556 VSS.n891 VSS.n888 585
R557 VSS.n2093 VSS.n2092 585
R558 VSS.n2094 VSS.n2093 585
R559 VSS.n2091 VSS.n892 585
R560 VSS.n892 VSS.n890 585
R561 VSS.n2090 VSS.n2089 585
R562 VSS.n2089 VSS.n2088 585
R563 VSS.n895 VSS.n894 585
R564 VSS.n2087 VSS.n895 585
R565 VSS.n2085 VSS.n2084 585
R566 VSS.n2086 VSS.n2085 585
R567 VSS.n2083 VSS.n900 585
R568 VSS.n900 VSS.n899 585
R569 VSS.n2554 VSS.n2553 585
R570 VSS.n2552 VSS.n100 585
R571 VSS.n2551 VSS.n99 585
R572 VSS.n2556 VSS.n99 585
R573 VSS.n2550 VSS.n2549 585
R574 VSS.n2548 VSS.n2547 585
R575 VSS.n2546 VSS.n2545 585
R576 VSS.n2544 VSS.n2543 585
R577 VSS.n2542 VSS.n2541 585
R578 VSS.n2540 VSS.n2539 585
R579 VSS.n2538 VSS.n2537 585
R580 VSS.n2536 VSS.n2535 585
R581 VSS.n2534 VSS.n2533 585
R582 VSS.n2532 VSS.n2531 585
R583 VSS.n2530 VSS.n2529 585
R584 VSS.n2528 VSS.n2527 585
R585 VSS.n2526 VSS.n2525 585
R586 VSS.n2518 VSS.n2500 585
R587 VSS.n2520 VSS.n2519 585
R588 VSS.n2517 VSS.n2516 585
R589 VSS.n2515 VSS.n2514 585
R590 VSS.n2504 VSS.n2503 585
R591 VSS.n2506 VSS.n2505 585
R592 VSS.n2509 VSS.n2508 585
R593 VSS.n79 VSS.n76 585
R594 VSS.n2559 VSS.n2558 585
R595 VSS.n78 VSS.n77 585
R596 VSS.n2467 VSS.n2466 585
R597 VSS.n2469 VSS.n2468 585
R598 VSS.n2471 VSS.n2470 585
R599 VSS.n2473 VSS.n2472 585
R600 VSS.n2475 VSS.n2474 585
R601 VSS.n2477 VSS.n2476 585
R602 VSS.n2479 VSS.n2478 585
R603 VSS.n2481 VSS.n2480 585
R604 VSS.n2483 VSS.n2482 585
R605 VSS.n2485 VSS.n2484 585
R606 VSS.n2487 VSS.n2486 585
R607 VSS.n2489 VSS.n2488 585
R608 VSS.n2491 VSS.n2490 585
R609 VSS.n2492 VSS.n106 585
R610 VSS.n106 VSS.n80 585
R611 VSS.n2494 VSS.n2493 585
R612 VSS.n2495 VSS.n2494 585
R613 VSS.n2465 VSS.n105 585
R614 VSS.n105 VSS.n104 585
R615 VSS.n2464 VSS.n2463 585
R616 VSS.n2463 VSS.n2462 585
R617 VSS.n108 VSS.n107 585
R618 VSS.n109 VSS.n108 585
R619 VSS.n2455 VSS.n2454 585
R620 VSS.n2456 VSS.n2455 585
R621 VSS.n2453 VSS.n113 585
R622 VSS.n117 VSS.n113 585
R623 VSS.n2452 VSS.n2451 585
R624 VSS.n2451 VSS.n2450 585
R625 VSS.n115 VSS.n114 585
R626 VSS.n116 VSS.n115 585
R627 VSS.n2443 VSS.n2442 585
R628 VSS.n2444 VSS.n2443 585
R629 VSS.n2441 VSS.n121 585
R630 VSS.n125 VSS.n121 585
R631 VSS.n2440 VSS.n2439 585
R632 VSS.n2439 VSS.n2438 585
R633 VSS.n123 VSS.n122 585
R634 VSS.n124 VSS.n123 585
R635 VSS.n2431 VSS.n2430 585
R636 VSS.n2432 VSS.n2431 585
R637 VSS.n2429 VSS.n129 585
R638 VSS.n133 VSS.n129 585
R639 VSS.n2428 VSS.n2427 585
R640 VSS.n2427 VSS.n2426 585
R641 VSS.n131 VSS.n130 585
R642 VSS.n132 VSS.n131 585
R643 VSS.n2419 VSS.n2418 585
R644 VSS.n2420 VSS.n2419 585
R645 VSS.n2417 VSS.n137 585
R646 VSS.n141 VSS.n137 585
R647 VSS.n2416 VSS.n2415 585
R648 VSS.n2415 VSS.n2414 585
R649 VSS.n139 VSS.n138 585
R650 VSS.n140 VSS.n139 585
R651 VSS.n2407 VSS.n2406 585
R652 VSS.n2408 VSS.n2407 585
R653 VSS.n2405 VSS.n145 585
R654 VSS.n149 VSS.n145 585
R655 VSS.n2404 VSS.n2403 585
R656 VSS.n2403 VSS.n2402 585
R657 VSS.n147 VSS.n146 585
R658 VSS.n148 VSS.n147 585
R659 VSS.n2395 VSS.n2394 585
R660 VSS.n2396 VSS.n2395 585
R661 VSS.n2393 VSS.n154 585
R662 VSS.n154 VSS.n153 585
R663 VSS.n2392 VSS.n2391 585
R664 VSS.n2391 VSS.n2390 585
R665 VSS.n156 VSS.n155 585
R666 VSS.n157 VSS.n156 585
R667 VSS.n2383 VSS.n2382 585
R668 VSS.n2384 VSS.n2383 585
R669 VSS.n2381 VSS.n162 585
R670 VSS.n162 VSS.n161 585
R671 VSS.n2380 VSS.n2379 585
R672 VSS.n2379 VSS.n2378 585
R673 VSS.n164 VSS.n163 585
R674 VSS.n165 VSS.n164 585
R675 VSS.n2371 VSS.n2370 585
R676 VSS.n2372 VSS.n2371 585
R677 VSS.n2369 VSS.n170 585
R678 VSS.n170 VSS.n169 585
R679 VSS.n2368 VSS.n2367 585
R680 VSS.n2367 VSS.n2366 585
R681 VSS.n172 VSS.n171 585
R682 VSS.n173 VSS.n172 585
R683 VSS.n2359 VSS.n2358 585
R684 VSS.n2360 VSS.n2359 585
R685 VSS.n2357 VSS.n178 585
R686 VSS.n178 VSS.n177 585
R687 VSS.n2356 VSS.n2355 585
R688 VSS.n2355 VSS.n2354 585
R689 VSS.n180 VSS.n179 585
R690 VSS.n2347 VSS.n180 585
R691 VSS.n2346 VSS.n2345 585
R692 VSS.n2348 VSS.n2346 585
R693 VSS.n2344 VSS.n185 585
R694 VSS.n185 VSS.n184 585
R695 VSS.n2343 VSS.n2342 585
R696 VSS.n2342 VSS.n2341 585
R697 VSS.n187 VSS.n186 585
R698 VSS.n2334 VSS.n187 585
R699 VSS.n2333 VSS.n2332 585
R700 VSS.n2335 VSS.n2333 585
R701 VSS.n2331 VSS.n192 585
R702 VSS.n192 VSS.n191 585
R703 VSS.n2330 VSS.n2329 585
R704 VSS.n2329 VSS.n2328 585
R705 VSS.n194 VSS.n193 585
R706 VSS.n2321 VSS.n194 585
R707 VSS.n2320 VSS.n2319 585
R708 VSS.n2322 VSS.n2320 585
R709 VSS.n2318 VSS.n199 585
R710 VSS.n199 VSS.n198 585
R711 VSS.n2317 VSS.n2316 585
R712 VSS.n2316 VSS.n2315 585
R713 VSS.n201 VSS.n200 585
R714 VSS.n2308 VSS.n201 585
R715 VSS.n2307 VSS.n2306 585
R716 VSS.n2309 VSS.n2307 585
R717 VSS.n2305 VSS.n206 585
R718 VSS.n206 VSS.n205 585
R719 VSS.n2304 VSS.n2303 585
R720 VSS.n2303 VSS.n2302 585
R721 VSS.n208 VSS.n207 585
R722 VSS.n2294 VSS.n208 585
R723 VSS.n442 VSS.n441 585
R724 VSS.n2296 VSS.n442 585
R725 VSS.n440 VSS.n213 585
R726 VSS.n213 VSS.n212 585
R727 VSS.n439 VSS.n438 585
R728 VSS.n438 VSS.n437 585
R729 VSS.n215 VSS.n214 585
R730 VSS.n216 VSS.n215 585
R731 VSS.n430 VSS.n429 585
R732 VSS.n431 VSS.n430 585
R733 VSS.n428 VSS.n221 585
R734 VSS.n427 VSS.n426 585
R735 VSS.n424 VSS.n222 585
R736 VSS.n422 VSS.n421 585
R737 VSS.n420 VSS.n223 585
R738 VSS.n419 VSS.n418 585
R739 VSS.n416 VSS.n224 585
R740 VSS.n414 VSS.n413 585
R741 VSS.n412 VSS.n225 585
R742 VSS.n411 VSS.n410 585
R743 VSS.n408 VSS.n226 585
R744 VSS.n406 VSS.n405 585
R745 VSS.n404 VSS.n227 585
R746 VSS.n403 VSS.n402 585
R747 VSS.n400 VSS.n228 585
R748 VSS.n398 VSS.n397 585
R749 VSS.n230 VSS.n229 585
R750 VSS.n292 VSS.n291 585
R751 VSS.n289 VSS.n232 585
R752 VSS.n287 VSS.n286 585
R753 VSS.n234 VSS.n233 585
R754 VSS.n280 VSS.n279 585
R755 VSS.n277 VSS.n236 585
R756 VSS.n275 VSS.n274 585
R757 VSS.n271 VSS.n237 585
R758 VSS.n270 VSS.n269 585
R759 VSS.n267 VSS.n238 585
R760 VSS.n265 VSS.n264 585
R761 VSS.n263 VSS.n239 585
R762 VSS.n262 VSS.n261 585
R763 VSS.n259 VSS.n240 585
R764 VSS.n257 VSS.n256 585
R765 VSS.n255 VSS.n241 585
R766 VSS.n254 VSS.n253 585
R767 VSS.n251 VSS.n242 585
R768 VSS.n249 VSS.n248 585
R769 VSS.n247 VSS.n243 585
R770 VSS.n246 VSS.n245 585
R771 VSS.n219 VSS.n218 585
R772 VSS.n220 VSS.n219 585
R773 VSS.n433 VSS.n432 585
R774 VSS.n432 VSS.n431 585
R775 VSS.n434 VSS.n217 585
R776 VSS.n217 VSS.n216 585
R777 VSS.n436 VSS.n435 585
R778 VSS.n437 VSS.n436 585
R779 VSS.n211 VSS.n210 585
R780 VSS.n212 VSS.n211 585
R781 VSS.n2298 VSS.n2297 585
R782 VSS.n2297 VSS.n2296 585
R783 VSS.n2299 VSS.n209 585
R784 VSS.n2294 VSS.n209 585
R785 VSS.n2301 VSS.n2300 585
R786 VSS.n2302 VSS.n2301 585
R787 VSS.n204 VSS.n203 585
R788 VSS.n205 VSS.n204 585
R789 VSS.n2311 VSS.n2310 585
R790 VSS.n2310 VSS.n2309 585
R791 VSS.n2312 VSS.n202 585
R792 VSS.n2308 VSS.n202 585
R793 VSS.n2314 VSS.n2313 585
R794 VSS.n2315 VSS.n2314 585
R795 VSS.n197 VSS.n196 585
R796 VSS.n198 VSS.n197 585
R797 VSS.n2324 VSS.n2323 585
R798 VSS.n2323 VSS.n2322 585
R799 VSS.n2325 VSS.n195 585
R800 VSS.n2321 VSS.n195 585
R801 VSS.n2327 VSS.n2326 585
R802 VSS.n2328 VSS.n2327 585
R803 VSS.n190 VSS.n189 585
R804 VSS.n191 VSS.n190 585
R805 VSS.n2337 VSS.n2336 585
R806 VSS.n2336 VSS.n2335 585
R807 VSS.n2338 VSS.n188 585
R808 VSS.n2334 VSS.n188 585
R809 VSS.n2340 VSS.n2339 585
R810 VSS.n2341 VSS.n2340 585
R811 VSS.n183 VSS.n182 585
R812 VSS.n184 VSS.n183 585
R813 VSS.n2350 VSS.n2349 585
R814 VSS.n2349 VSS.n2348 585
R815 VSS.n2351 VSS.n181 585
R816 VSS.n2347 VSS.n181 585
R817 VSS.n2353 VSS.n2352 585
R818 VSS.n2354 VSS.n2353 585
R819 VSS.n176 VSS.n175 585
R820 VSS.n177 VSS.n176 585
R821 VSS.n2362 VSS.n2361 585
R822 VSS.n2361 VSS.n2360 585
R823 VSS.n2363 VSS.n174 585
R824 VSS.n174 VSS.n173 585
R825 VSS.n2365 VSS.n2364 585
R826 VSS.n2366 VSS.n2365 585
R827 VSS.n168 VSS.n167 585
R828 VSS.n169 VSS.n168 585
R829 VSS.n2374 VSS.n2373 585
R830 VSS.n2373 VSS.n2372 585
R831 VSS.n2375 VSS.n166 585
R832 VSS.n166 VSS.n165 585
R833 VSS.n2377 VSS.n2376 585
R834 VSS.n2378 VSS.n2377 585
R835 VSS.n160 VSS.n159 585
R836 VSS.n161 VSS.n160 585
R837 VSS.n2386 VSS.n2385 585
R838 VSS.n2385 VSS.n2384 585
R839 VSS.n2387 VSS.n158 585
R840 VSS.n158 VSS.n157 585
R841 VSS.n2389 VSS.n2388 585
R842 VSS.n2390 VSS.n2389 585
R843 VSS.n152 VSS.n151 585
R844 VSS.n153 VSS.n152 585
R845 VSS.n2398 VSS.n2397 585
R846 VSS.n2397 VSS.n2396 585
R847 VSS.n2399 VSS.n150 585
R848 VSS.n150 VSS.n148 585
R849 VSS.n2401 VSS.n2400 585
R850 VSS.n2402 VSS.n2401 585
R851 VSS.n144 VSS.n143 585
R852 VSS.n149 VSS.n144 585
R853 VSS.n2410 VSS.n2409 585
R854 VSS.n2409 VSS.n2408 585
R855 VSS.n2411 VSS.n142 585
R856 VSS.n142 VSS.n140 585
R857 VSS.n2413 VSS.n2412 585
R858 VSS.n2414 VSS.n2413 585
R859 VSS.n136 VSS.n135 585
R860 VSS.n141 VSS.n136 585
R861 VSS.n2422 VSS.n2421 585
R862 VSS.n2421 VSS.n2420 585
R863 VSS.n2423 VSS.n134 585
R864 VSS.n134 VSS.n132 585
R865 VSS.n2425 VSS.n2424 585
R866 VSS.n2426 VSS.n2425 585
R867 VSS.n128 VSS.n127 585
R868 VSS.n133 VSS.n128 585
R869 VSS.n2434 VSS.n2433 585
R870 VSS.n2433 VSS.n2432 585
R871 VSS.n2435 VSS.n126 585
R872 VSS.n126 VSS.n124 585
R873 VSS.n2437 VSS.n2436 585
R874 VSS.n2438 VSS.n2437 585
R875 VSS.n120 VSS.n119 585
R876 VSS.n125 VSS.n120 585
R877 VSS.n2446 VSS.n2445 585
R878 VSS.n2445 VSS.n2444 585
R879 VSS.n2447 VSS.n118 585
R880 VSS.n118 VSS.n116 585
R881 VSS.n2449 VSS.n2448 585
R882 VSS.n2450 VSS.n2449 585
R883 VSS.n112 VSS.n111 585
R884 VSS.n117 VSS.n112 585
R885 VSS.n2458 VSS.n2457 585
R886 VSS.n2457 VSS.n2456 585
R887 VSS.n2459 VSS.n110 585
R888 VSS.n110 VSS.n109 585
R889 VSS.n2461 VSS.n2460 585
R890 VSS.n2462 VSS.n2461 585
R891 VSS.n103 VSS.n102 585
R892 VSS.n104 VSS.n103 585
R893 VSS.n2497 VSS.n2496 585
R894 VSS.n2496 VSS.n2495 585
R895 VSS.n2498 VSS.n101 585
R896 VSS.n101 VSS.n80 585
R897 VSS.n1134 VSS.n1133 585
R898 VSS.n1131 VSS.n953 585
R899 VSS.n1130 VSS.n1129 585
R900 VSS.n1130 VSS.n890 585
R901 VSS.n1128 VSS.n954 585
R902 VSS.n1127 VSS.n1126 585
R903 VSS.n1124 VSS.n955 585
R904 VSS.n1122 VSS.n1121 585
R905 VSS.n1120 VSS.n956 585
R906 VSS.n1119 VSS.n1118 585
R907 VSS.n1116 VSS.n957 585
R908 VSS.n1114 VSS.n1113 585
R909 VSS.n1112 VSS.n958 585
R910 VSS.n1111 VSS.n1110 585
R911 VSS.n1108 VSS.n959 585
R912 VSS.n1106 VSS.n1105 585
R913 VSS.n1104 VSS.n960 585
R914 VSS.n1103 VSS.n1102 585
R915 VSS.n1100 VSS.n961 585
R916 VSS.n1098 VSS.n1097 585
R917 VSS.n1096 VSS.n962 585
R918 VSS.n1095 VSS.n1094 585
R919 VSS.n1092 VSS.n963 585
R920 VSS.n1090 VSS.n1089 585
R921 VSS.n1088 VSS.n964 585
R922 VSS.n1087 VSS.n1086 585
R923 VSS.n1084 VSS.n965 585
R924 VSS.n1082 VSS.n1081 585
R925 VSS.n1080 VSS.n966 585
R926 VSS.n1079 VSS.n1078 585
R927 VSS.n1076 VSS.n967 585
R928 VSS.n1074 VSS.n1073 585
R929 VSS.n1072 VSS.n968 585
R930 VSS.n1071 VSS.n1070 585
R931 VSS.n1068 VSS.n969 585
R932 VSS.n1066 VSS.n1065 585
R933 VSS.n1064 VSS.n970 585
R934 VSS.n1063 VSS.n1062 585
R935 VSS.n1060 VSS.n971 585
R936 VSS.n1058 VSS.n1057 585
R937 VSS.n1056 VSS.n972 585
R938 VSS.n1055 VSS.n1054 585
R939 VSS.n1052 VSS.n973 585
R940 VSS.n1050 VSS.n1049 585
R941 VSS.n1048 VSS.n974 585
R942 VSS.n1047 VSS.n1046 585
R943 VSS.n1044 VSS.n975 585
R944 VSS.n1042 VSS.n1041 585
R945 VSS.n1040 VSS.n976 585
R946 VSS.n1039 VSS.n1038 585
R947 VSS.n1036 VSS.n977 585
R948 VSS.n1034 VSS.n1033 585
R949 VSS.n1032 VSS.n978 585
R950 VSS.n1031 VSS.n1030 585
R951 VSS.n1028 VSS.n979 585
R952 VSS.n1026 VSS.n1025 585
R953 VSS.n1024 VSS.n980 585
R954 VSS.n1023 VSS.n1022 585
R955 VSS.n1020 VSS.n981 585
R956 VSS.n1018 VSS.n1017 585
R957 VSS.n1016 VSS.n982 585
R958 VSS.n1015 VSS.n1014 585
R959 VSS.n1012 VSS.n983 585
R960 VSS.n1010 VSS.n1009 585
R961 VSS.n1008 VSS.n984 585
R962 VSS.n1007 VSS.n1006 585
R963 VSS.n1004 VSS.n985 585
R964 VSS.n1002 VSS.n1001 585
R965 VSS.n1000 VSS.n986 585
R966 VSS.n999 VSS.n998 585
R967 VSS.n996 VSS.n987 585
R968 VSS.n994 VSS.n993 585
R969 VSS.n992 VSS.n988 585
R970 VSS.n991 VSS.n990 585
R971 VSS.n887 VSS.n886 585
R972 VSS.n890 VSS.n887 585
R973 VSS.n2097 VSS.n2096 585
R974 VSS.n2096 VSS.n2095 585
R975 VSS.n884 VSS.n882 585
R976 VSS.n2024 VSS.n882 585
R977 VSS.n2102 VSS.n2101 585
R978 VSS.n2103 VSS.n2102 585
R979 VSS.n883 VSS.n881 585
R980 VSS.n881 VSS.n879 585
R981 VSS.n870 VSS.n868 585
R982 VSS.n873 VSS.n870 585
R983 VSS.n2113 VSS.n2112 585
R984 VSS.n2112 VSS.n2111 585
R985 VSS.n869 VSS.n867 585
R986 VSS.n1957 VSS.n869 585
R987 VSS.n1958 VSS.n865 585
R988 VSS.n1959 VSS.n1958 585
R989 VSS.n2117 VSS.n863 585
R990 VSS.n863 VSS.n861 585
R991 VSS.n2119 VSS.n2118 585
R992 VSS.n2120 VSS.n2119 585
R993 VSS.n864 VSS.n862 585
R994 VSS.n862 VSS.n781 585
R995 VSS.n772 VSS.n771 585
R996 VSS.n775 VSS.n772 585
R997 VSS.n2131 VSS.n2130 585
R998 VSS.n2130 VSS.n2129 585
R999 VSS.n2132 VSS.n769 585
R1000 VSS.n1187 VSS.n769 585
R1001 VSS.n2134 VSS.n2133 585
R1002 VSS.n2135 VSS.n2134 585
R1003 VSS.n770 VSS.n768 585
R1004 VSS.n768 VSS.n765 585
R1005 VSS.n1891 VSS.n757 585
R1006 VSS.n759 VSS.n757 585
R1007 VSS.n2145 VSS.n2144 585
R1008 VSS.n2144 VSS.n2143 585
R1009 VSS.n2146 VSS.n753 585
R1010 VSS.n840 VSS.n753 585
R1011 VSS.n2148 VSS.n2147 585
R1012 VSS.n2149 VSS.n2148 585
R1013 VSS.n754 VSS.n752 585
R1014 VSS.n752 VSS.n749 585
R1015 VSS.n1903 VSS.n1902 585
R1016 VSS.n1904 VSS.n1903 585
R1017 VSS.n1325 VSS.n1324 585
R1018 VSS.n1324 VSS.n700 585
R1019 VSS.n1331 VSS.n1330 585
R1020 VSS.n1330 VSS.n1329 585
R1021 VSS.n1327 VSS.n1326 585
R1022 VSS.n1327 VSS.n694 585
R1023 VSS.n679 VSS.n678 585
R1024 VSS.n2163 VSS.n679 585
R1025 VSS.n2166 VSS.n2165 585
R1026 VSS.n2165 VSS.n2164 585
R1027 VSS.n2167 VSS.n676 585
R1028 VSS.n676 VSS.n674 585
R1029 VSS.n2169 VSS.n2168 585
R1030 VSS.n2170 VSS.n2169 585
R1031 VSS.n677 VSS.n675 585
R1032 VSS.n1409 VSS.n675 585
R1033 VSS.n1817 VSS.n1815 585
R1034 VSS.n1815 VSS.n1814 585
R1035 VSS.n1823 VSS.n1822 585
R1036 VSS.n1824 VSS.n1823 585
R1037 VSS.n1816 VSS.n1407 585
R1038 VSS.n1407 VSS.n1404 585
R1039 VSS.n1396 VSS.n1394 585
R1040 VSS.n1398 VSS.n1396 585
R1041 VSS.n1834 VSS.n1833 585
R1042 VSS.n1833 VSS.n1832 585
R1043 VSS.n1395 VSS.n1393 585
R1044 VSS.n1743 VSS.n1395 585
R1045 VSS.n1730 VSS.n1434 585
R1046 VSS.n1434 VSS.n1427 585
R1047 VSS.n1734 VSS.n1733 585
R1048 VSS.n1735 VSS.n1734 585
R1049 VSS.n1728 VSS.n1433 585
R1050 VSS.n1656 VSS.n1433 585
R1051 VSS.n1727 VSS.n1726 585
R1052 VSS.n1436 VSS.n1435 585
R1053 VSS.n1653 VSS.n1652 585
R1054 VSS.n1651 VSS.n1472 585
R1055 VSS.n1650 VSS.n1649 585
R1056 VSS.n1648 VSS.n1647 585
R1057 VSS.n1646 VSS.n1645 585
R1058 VSS.n1644 VSS.n1643 585
R1059 VSS.n1642 VSS.n1641 585
R1060 VSS.n1640 VSS.n1639 585
R1061 VSS.n1638 VSS.n1637 585
R1062 VSS.n1636 VSS.n1635 585
R1063 VSS.n1634 VSS.n1633 585
R1064 VSS.n1632 VSS.n1631 585
R1065 VSS.n1630 VSS.n1629 585
R1066 VSS.n1628 VSS.n1627 585
R1067 VSS.n1626 VSS.n1625 585
R1068 VSS.n1624 VSS.n1623 585
R1069 VSS.n1622 VSS.n1621 585
R1070 VSS.n1620 VSS.n1619 585
R1071 VSS.n1618 VSS.n1617 585
R1072 VSS.n1616 VSS.n1615 585
R1073 VSS.n1614 VSS.n1613 585
R1074 VSS.n1612 VSS.n1611 585
R1075 VSS.n1610 VSS.n1609 585
R1076 VSS.n1608 VSS.n1607 585
R1077 VSS.n1606 VSS.n1605 585
R1078 VSS.n1604 VSS.n1603 585
R1079 VSS.n1602 VSS.n1601 585
R1080 VSS.n1600 VSS.n1599 585
R1081 VSS.n1598 VSS.n1597 585
R1082 VSS.n1596 VSS.n1595 585
R1083 VSS.n1594 VSS.n1593 585
R1084 VSS.n1592 VSS.n1591 585
R1085 VSS.n1590 VSS.n1589 585
R1086 VSS.n1588 VSS.n1587 585
R1087 VSS.n1586 VSS.n1585 585
R1088 VSS.n1584 VSS.n1583 585
R1089 VSS.n1582 VSS.n1581 585
R1090 VSS.n1580 VSS.n1579 585
R1091 VSS.n1578 VSS.n1577 585
R1092 VSS.n1576 VSS.n1575 585
R1093 VSS.n1574 VSS.n1573 585
R1094 VSS.n1572 VSS.n1571 585
R1095 VSS.n1570 VSS.n1569 585
R1096 VSS.n1568 VSS.n1567 585
R1097 VSS.n1566 VSS.n1565 585
R1098 VSS.n1564 VSS.n1563 585
R1099 VSS.n1562 VSS.n1561 585
R1100 VSS.n1560 VSS.n1559 585
R1101 VSS.n1558 VSS.n1557 585
R1102 VSS.n1556 VSS.n1555 585
R1103 VSS.n1554 VSS.n1553 585
R1104 VSS.n1552 VSS.n1551 585
R1105 VSS.n1550 VSS.n1549 585
R1106 VSS.n1548 VSS.n1547 585
R1107 VSS.n1546 VSS.n1545 585
R1108 VSS.n1544 VSS.n1543 585
R1109 VSS.n1542 VSS.n1541 585
R1110 VSS.n1540 VSS.n1539 585
R1111 VSS.n1538 VSS.n1537 585
R1112 VSS.n1536 VSS.n1535 585
R1113 VSS.n1534 VSS.n1533 585
R1114 VSS.n1532 VSS.n1531 585
R1115 VSS.n1530 VSS.n1529 585
R1116 VSS.n1528 VSS.n1527 585
R1117 VSS.n1526 VSS.n1525 585
R1118 VSS.n1524 VSS.n1523 585
R1119 VSS.n1522 VSS.n1521 585
R1120 VSS.n1520 VSS.n1519 585
R1121 VSS.n1518 VSS.n1517 585
R1122 VSS.n1516 VSS.n1515 585
R1123 VSS.n1514 VSS.n1513 585
R1124 VSS.n1512 VSS.n1511 585
R1125 VSS.n2161 VSS.n2160 585
R1126 VSS.n2162 VSS.n2161 585
R1127 VSS.n697 VSS.n695 585
R1128 VSS.n705 VSS.n704 585
R1129 VSS.n707 VSS.n706 585
R1130 VSS.n709 VSS.n708 585
R1131 VSS.n711 VSS.n710 585
R1132 VSS.n713 VSS.n712 585
R1133 VSS.n715 VSS.n714 585
R1134 VSS.n717 VSS.n716 585
R1135 VSS.n719 VSS.n718 585
R1136 VSS.n721 VSS.n720 585
R1137 VSS.n723 VSS.n722 585
R1138 VSS.n725 VSS.n724 585
R1139 VSS.n727 VSS.n726 585
R1140 VSS.n729 VSS.n728 585
R1141 VSS.n731 VSS.n730 585
R1142 VSS.n733 VSS.n732 585
R1143 VSS.n735 VSS.n734 585
R1144 VSS.n737 VSS.n736 585
R1145 VSS.n739 VSS.n738 585
R1146 VSS.n741 VSS.n740 585
R1147 VSS.n743 VSS.n742 585
R1148 VSS.n745 VSS.n744 585
R1149 VSS.n746 VSS.n702 585
R1150 VSS.n1328 VSS.n702 585
R1151 VSS.n2155 VSS.n2154 585
R1152 VSS.n2156 VSS.n2155 585
R1153 VSS.n2153 VSS.n703 585
R1154 VSS.n1905 VSS.n703 585
R1155 VSS.n2152 VSS.n2151 585
R1156 VSS.n2151 VSS.n2150 585
R1157 VSS.n748 VSS.n747 585
R1158 VSS.n751 VSS.n748 585
R1159 VSS.n762 VSS.n760 585
R1160 VSS.n841 VSS.n760 585
R1161 VSS.n2141 VSS.n2140 585
R1162 VSS.n2142 VSS.n2141 585
R1163 VSS.n2139 VSS.n761 585
R1164 VSS.n829 VSS.n761 585
R1165 VSS.n2138 VSS.n2137 585
R1166 VSS.n2137 VSS.n2136 585
R1167 VSS.n764 VSS.n763 585
R1168 VSS.n767 VSS.n764 585
R1169 VSS.n778 VSS.n776 585
R1170 VSS.n776 VSS.n773 585
R1171 VSS.n2127 VSS.n2126 585
R1172 VSS.n2128 VSS.n2127 585
R1173 VSS.n2125 VSS.n777 585
R1174 VSS.n2124 VSS.n2123 585
R1175 VSS.n780 VSS.n779 585
R1176 VSS.n2121 VSS.n780 585
R1177 VSS.n793 VSS.n792 585
R1178 VSS.n795 VSS.n794 585
R1179 VSS.n797 VSS.n796 585
R1180 VSS.n799 VSS.n798 585
R1181 VSS.n801 VSS.n800 585
R1182 VSS.n803 VSS.n802 585
R1183 VSS.n805 VSS.n804 585
R1184 VSS.n807 VSS.n806 585
R1185 VSS.n809 VSS.n808 585
R1186 VSS.n811 VSS.n810 585
R1187 VSS.n813 VSS.n812 585
R1188 VSS.n815 VSS.n814 585
R1189 VSS.n817 VSS.n816 585
R1190 VSS.n819 VSS.n818 585
R1191 VSS.n821 VSS.n820 585
R1192 VSS.n823 VSS.n822 585
R1193 VSS.n825 VSS.n824 585
R1194 VSS.n827 VSS.n826 585
R1195 VSS.n828 VSS.n791 585
R1196 VSS.n857 VSS.n856 585
R1197 VSS.n855 VSS.n774 585
R1198 VSS.n2128 VSS.n774 585
R1199 VSS.n854 VSS.n853 585
R1200 VSS.n853 VSS.n773 585
R1201 VSS.n852 VSS.n851 585
R1202 VSS.n852 VSS.n767 585
R1203 VSS.n849 VSS.n766 585
R1204 VSS.n2136 VSS.n766 585
R1205 VSS.n831 VSS.n830 585
R1206 VSS.n830 VSS.n829 585
R1207 VSS.n844 VSS.n758 585
R1208 VSS.n2142 VSS.n758 585
R1209 VSS.n843 VSS.n842 585
R1210 VSS.n842 VSS.n841 585
R1211 VSS.n839 VSS.n838 585
R1212 VSS.n839 VSS.n751 585
R1213 VSS.n837 VSS.n750 585
R1214 VSS.n2150 VSS.n750 585
R1215 VSS.n834 VSS.n699 585
R1216 VSS.n1905 VSS.n699 585
R1217 VSS.n2158 VSS.n2157 585
R1218 VSS.n2157 VSS.n2156 585
R1219 VSS.n2159 VSS.n696 585
R1220 VSS.n1328 VSS.n696 585
R1221 VSS.n432 VSS.n217 394
R1222 VSS.n436 VSS.n217 394
R1223 VSS.n436 VSS.n211 394
R1224 VSS.n2297 VSS.n211 394
R1225 VSS.n2297 VSS.n209 394
R1226 VSS.n2301 VSS.n209 394
R1227 VSS.n2301 VSS.n204 394
R1228 VSS.n2310 VSS.n204 394
R1229 VSS.n2310 VSS.n202 394
R1230 VSS.n2314 VSS.n202 394
R1231 VSS.n2314 VSS.n197 394
R1232 VSS.n2323 VSS.n197 394
R1233 VSS.n2323 VSS.n195 394
R1234 VSS.n2327 VSS.n195 394
R1235 VSS.n2327 VSS.n190 394
R1236 VSS.n2336 VSS.n190 394
R1237 VSS.n2336 VSS.n188 394
R1238 VSS.n2340 VSS.n188 394
R1239 VSS.n2340 VSS.n183 394
R1240 VSS.n2349 VSS.n183 394
R1241 VSS.n2349 VSS.n181 394
R1242 VSS.n2353 VSS.n181 394
R1243 VSS.n2353 VSS.n176 394
R1244 VSS.n2361 VSS.n176 394
R1245 VSS.n2361 VSS.n174 394
R1246 VSS.n2365 VSS.n174 394
R1247 VSS.n2365 VSS.n168 394
R1248 VSS.n2373 VSS.n168 394
R1249 VSS.n2373 VSS.n166 394
R1250 VSS.n2377 VSS.n166 394
R1251 VSS.n2377 VSS.n160 394
R1252 VSS.n2385 VSS.n160 394
R1253 VSS.n2385 VSS.n158 394
R1254 VSS.n2389 VSS.n158 394
R1255 VSS.n2389 VSS.n152 394
R1256 VSS.n2397 VSS.n152 394
R1257 VSS.n2397 VSS.n150 394
R1258 VSS.n2401 VSS.n150 394
R1259 VSS.n2401 VSS.n144 394
R1260 VSS.n2409 VSS.n144 394
R1261 VSS.n2409 VSS.n142 394
R1262 VSS.n2413 VSS.n142 394
R1263 VSS.n2413 VSS.n136 394
R1264 VSS.n2421 VSS.n136 394
R1265 VSS.n2421 VSS.n134 394
R1266 VSS.n2425 VSS.n134 394
R1267 VSS.n2425 VSS.n128 394
R1268 VSS.n2433 VSS.n128 394
R1269 VSS.n2433 VSS.n126 394
R1270 VSS.n2437 VSS.n126 394
R1271 VSS.n2437 VSS.n120 394
R1272 VSS.n2445 VSS.n120 394
R1273 VSS.n2445 VSS.n118 394
R1274 VSS.n2449 VSS.n118 394
R1275 VSS.n2449 VSS.n112 394
R1276 VSS.n2457 VSS.n112 394
R1277 VSS.n2457 VSS.n110 394
R1278 VSS.n2461 VSS.n110 394
R1279 VSS.n2461 VSS.n103 394
R1280 VSS.n2496 VSS.n103 394
R1281 VSS.n2496 VSS.n101 394
R1282 VSS.n245 VSS.n219 394
R1283 VSS.n249 VSS.n243 394
R1284 VSS.n253 VSS.n251 394
R1285 VSS.n257 VSS.n241 394
R1286 VSS.n261 VSS.n259 394
R1287 VSS.n265 VSS.n239 394
R1288 VSS.n269 VSS.n267 394
R1289 VSS.n275 VSS.n237 394
R1290 VSS.n279 VSS.n277 394
R1291 VSS.n287 VSS.n233 394
R1292 VSS.n291 VSS.n289 394
R1293 VSS.n398 VSS.n229 394
R1294 VSS.n402 VSS.n400 394
R1295 VSS.n406 VSS.n227 394
R1296 VSS.n410 VSS.n408 394
R1297 VSS.n414 VSS.n225 394
R1298 VSS.n418 VSS.n416 394
R1299 VSS.n422 VSS.n223 394
R1300 VSS.n426 VSS.n424 394
R1301 VSS.n430 VSS.n215 394
R1302 VSS.n438 VSS.n215 394
R1303 VSS.n438 VSS.n213 394
R1304 VSS.n442 VSS.n213 394
R1305 VSS.n442 VSS.n208 394
R1306 VSS.n2303 VSS.n208 394
R1307 VSS.n2303 VSS.n206 394
R1308 VSS.n2307 VSS.n206 394
R1309 VSS.n2307 VSS.n201 394
R1310 VSS.n2316 VSS.n201 394
R1311 VSS.n2316 VSS.n199 394
R1312 VSS.n2320 VSS.n199 394
R1313 VSS.n2320 VSS.n194 394
R1314 VSS.n2329 VSS.n194 394
R1315 VSS.n2329 VSS.n192 394
R1316 VSS.n2333 VSS.n192 394
R1317 VSS.n2333 VSS.n187 394
R1318 VSS.n2342 VSS.n187 394
R1319 VSS.n2342 VSS.n185 394
R1320 VSS.n2346 VSS.n185 394
R1321 VSS.n2346 VSS.n180 394
R1322 VSS.n2355 VSS.n180 394
R1323 VSS.n2355 VSS.n178 394
R1324 VSS.n2359 VSS.n178 394
R1325 VSS.n2359 VSS.n172 394
R1326 VSS.n2367 VSS.n172 394
R1327 VSS.n2367 VSS.n170 394
R1328 VSS.n2371 VSS.n170 394
R1329 VSS.n2371 VSS.n164 394
R1330 VSS.n2379 VSS.n164 394
R1331 VSS.n2379 VSS.n162 394
R1332 VSS.n2383 VSS.n162 394
R1333 VSS.n2383 VSS.n156 394
R1334 VSS.n2391 VSS.n156 394
R1335 VSS.n2391 VSS.n154 394
R1336 VSS.n2395 VSS.n154 394
R1337 VSS.n2395 VSS.n147 394
R1338 VSS.n2403 VSS.n147 394
R1339 VSS.n2403 VSS.n145 394
R1340 VSS.n2407 VSS.n145 394
R1341 VSS.n2407 VSS.n139 394
R1342 VSS.n2415 VSS.n139 394
R1343 VSS.n2415 VSS.n137 394
R1344 VSS.n2419 VSS.n137 394
R1345 VSS.n2419 VSS.n131 394
R1346 VSS.n2427 VSS.n131 394
R1347 VSS.n2427 VSS.n129 394
R1348 VSS.n2431 VSS.n129 394
R1349 VSS.n2431 VSS.n123 394
R1350 VSS.n2439 VSS.n123 394
R1351 VSS.n2439 VSS.n121 394
R1352 VSS.n2443 VSS.n121 394
R1353 VSS.n2443 VSS.n115 394
R1354 VSS.n2451 VSS.n115 394
R1355 VSS.n2451 VSS.n113 394
R1356 VSS.n2455 VSS.n113 394
R1357 VSS.n2455 VSS.n108 394
R1358 VSS.n2463 VSS.n108 394
R1359 VSS.n2463 VSS.n105 394
R1360 VSS.n2494 VSS.n105 394
R1361 VSS.n2494 VSS.n106 394
R1362 VSS.n100 VSS.n99 394
R1363 VSS.n2549 VSS.n99 394
R1364 VSS.n2547 VSS.n2546 394
R1365 VSS.n2543 VSS.n2542 394
R1366 VSS.n2539 VSS.n2538 394
R1367 VSS.n2535 VSS.n2534 394
R1368 VSS.n2531 VSS.n2530 394
R1369 VSS.n2527 VSS.n2526 394
R1370 VSS.n2519 VSS.n2518 394
R1371 VSS.n2516 VSS.n2515 394
R1372 VSS.n2505 VSS.n2504 394
R1373 VSS.n2508 VSS.n79 394
R1374 VSS.n2558 VSS.n78 394
R1375 VSS.n2468 VSS.n2467 394
R1376 VSS.n2472 VSS.n2471 394
R1377 VSS.n2476 VSS.n2475 394
R1378 VSS.n2480 VSS.n2479 394
R1379 VSS.n2484 VSS.n2483 394
R1380 VSS.n2488 VSS.n2487 394
R1381 VSS.n2109 VSS.n874 394
R1382 VSS.n2109 VSS.n875 394
R1383 VSS.n2105 VSS.n875 394
R1384 VSS.n2105 VSS.n878 394
R1385 VSS.n891 VSS.n878 394
R1386 VSS.n2093 VSS.n891 394
R1387 VSS.n2093 VSS.n892 394
R1388 VSS.n2089 VSS.n892 394
R1389 VSS.n2089 VSS.n895 394
R1390 VSS.n2085 VSS.n895 394
R1391 VSS.n2085 VSS.n900 394
R1392 VSS.n2012 VSS.n1970 394
R1393 VSS.n2008 VSS.n2007 394
R1394 VSS.n2004 VSS.n2003 394
R1395 VSS.n2000 VSS.n1999 394
R1396 VSS.n1996 VSS.n1995 394
R1397 VSS.n1992 VSS.n1991 394
R1398 VSS.n1988 VSS.n1987 394
R1399 VSS.n1984 VSS.n1983 394
R1400 VSS.n1980 VSS.n1979 394
R1401 VSS.n1976 VSS.n1975 394
R1402 VSS.n1972 VSS.n925 394
R1403 VSS.n2016 VSS.n872 394
R1404 VSS.n2020 VSS.n872 394
R1405 VSS.n2020 VSS.n880 394
R1406 VSS.n2026 VSS.n880 394
R1407 VSS.n2027 VSS.n2026 394
R1408 VSS.n2027 VSS.n889 394
R1409 VSS.n2030 VSS.n889 394
R1410 VSS.n2030 VSS.n896 394
R1411 VSS.n897 VSS.n896 394
R1412 VSS.n898 VSS.n897 394
R1413 VSS.n2036 VSS.n898 394
R1414 VSS.n2078 VSS.n902 394
R1415 VSS.n2078 VSS.n913 394
R1416 VSS.n2074 VSS.n2073 394
R1417 VSS.n2070 VSS.n2069 394
R1418 VSS.n919 VSS.n918 394
R1419 VSS.n2062 VSS.n2061 394
R1420 VSS.n2058 VSS.n2057 394
R1421 VSS.n2053 VSS.n2052 394
R1422 VSS.n2049 VSS.n2048 394
R1423 VSS.n2045 VSS.n2044 394
R1424 VSS.n2041 VSS.n2040 394
R1425 VSS.n1722 VSS.n1430 394
R1426 VSS.n1737 VSS.n1430 394
R1427 VSS.n1737 VSS.n1428 394
R1428 VSS.n1741 VSS.n1428 394
R1429 VSS.n1741 VSS.n1399 394
R1430 VSS.n1830 VSS.n1399 394
R1431 VSS.n1830 VSS.n1400 394
R1432 VSS.n1826 VSS.n1400 394
R1433 VSS.n1826 VSS.n1403 394
R1434 VSS.n1812 VSS.n1403 394
R1435 VSS.n1812 VSS.n1410 394
R1436 VSS.n1718 VSS.n1658 394
R1437 VSS.n1716 VSS.n1715 394
R1438 VSS.n1713 VSS.n1661 394
R1439 VSS.n1709 VSS.n1708 394
R1440 VSS.n1706 VSS.n1664 394
R1441 VSS.n1702 VSS.n1701 394
R1442 VSS.n1699 VSS.n1667 394
R1443 VSS.n1695 VSS.n1694 394
R1444 VSS.n1692 VSS.n1670 394
R1445 VSS.n1688 VSS.n1687 394
R1446 VSS.n1685 VSS.n1673 394
R1447 VSS.n1677 VSS.n1655 394
R1448 VSS.n1677 VSS.n1431 394
R1449 VSS.n1674 VSS.n1431 394
R1450 VSS.n1674 VSS.n1426 394
R1451 VSS.n1745 VSS.n1426 394
R1452 VSS.n1745 VSS.n1397 394
R1453 VSS.n1752 VSS.n1397 394
R1454 VSS.n1752 VSS.n1405 394
R1455 VSS.n1758 VSS.n1405 394
R1456 VSS.n1758 VSS.n1408 394
R1457 VSS.n1422 VSS.n1408 394
R1458 VSS.n1806 VSS.n1805 394
R1459 VSS.n1805 VSS.n1412 394
R1460 VSS.n1801 VSS.n1799 394
R1461 VSS.n1797 VSS.n1414 394
R1462 VSS.n1793 VSS.n1791 394
R1463 VSS.n1789 VSS.n1416 394
R1464 VSS.n1785 VSS.n1783 394
R1465 VSS.n1781 VSS.n1418 394
R1466 VSS.n1777 VSS.n1775 394
R1467 VSS.n1773 VSS.n1420 394
R1468 VSS.n1769 VSS.n1767 394
R1469 VSS.n2190 VSS.n656 394
R1470 VSS.n2184 VSS.n656 394
R1471 VSS.n2184 VSS.n661 394
R1472 VSS.n2180 VSS.n661 394
R1473 VSS.n2180 VSS.n663 394
R1474 VSS.n1749 VSS.n663 394
R1475 VSS.n1749 VSS.n669 394
R1476 VSS.n2173 VSS.n669 394
R1477 VSS.n2173 VSS.n670 394
R1478 VSS.n1303 VSS.n670 394
R1479 VSS.n1306 VSS.n1303 394
R1480 VSS.n1309 VSS.n1306 394
R1481 VSS.n1310 VSS.n1309 394
R1482 VSS.n1310 VSS.n1301 394
R1483 VSS.n1314 VSS.n1301 394
R1484 VSS.n1317 VSS.n1314 394
R1485 VSS.n1907 VSS.n1317 394
R1486 VSS.n1907 VSS.n1318 394
R1487 VSS.n1321 VSS.n1318 394
R1488 VSS.n1321 VSS.n1191 394
R1489 VSS.n1920 VSS.n1191 394
R1490 VSS.n1920 VSS.n1190 394
R1491 VSS.n1925 VSS.n1190 394
R1492 VSS.n1925 VSS.n1188 394
R1493 VSS.n1929 VSS.n1188 394
R1494 VSS.n1929 VSS.n1186 394
R1495 VSS.n1933 VSS.n1186 394
R1496 VSS.n1933 VSS.n1184 394
R1497 VSS.n1937 VSS.n1184 394
R1498 VSS.n1938 VSS.n1937 394
R1499 VSS.n1941 VSS.n1938 394
R1500 VSS.n1941 VSS.n928 394
R1501 VSS.n1955 VSS.n928 394
R1502 VSS.n1955 VSS.n929 394
R1503 VSS.n936 VSS.n929 394
R1504 VSS.n939 VSS.n936 394
R1505 VSS.n1176 VSS.n939 394
R1506 VSS.n1176 VSS.n940 394
R1507 VSS.n1475 VSS.n1474 394
R1508 VSS.n1479 VSS.n1478 394
R1509 VSS.n1483 VSS.n1482 394
R1510 VSS.n1487 VSS.n1486 394
R1511 VSS.n1491 VSS.n1490 394
R1512 VSS.n1495 VSS.n1494 394
R1513 VSS.n1499 VSS.n1498 394
R1514 VSS.n1503 VSS.n1502 394
R1515 VSS.n1507 VSS.n1506 394
R1516 VSS.n1511 VSS.n1510 394
R1517 VSS.n1515 VSS.n1514 394
R1518 VSS.n1519 VSS.n1518 394
R1519 VSS.n1523 VSS.n1522 394
R1520 VSS.n1527 VSS.n1526 394
R1521 VSS.n1531 VSS.n1530 394
R1522 VSS.n1535 VSS.n1534 394
R1523 VSS.n1539 VSS.n1538 394
R1524 VSS.n1543 VSS.n1542 394
R1525 VSS.n1547 VSS.n1546 394
R1526 VSS.n1551 VSS.n1550 394
R1527 VSS.n1555 VSS.n1554 394
R1528 VSS.n1559 VSS.n1558 394
R1529 VSS.n1563 VSS.n1562 394
R1530 VSS.n1567 VSS.n1566 394
R1531 VSS.n1571 VSS.n1570 394
R1532 VSS.n1575 VSS.n1574 394
R1533 VSS.n1579 VSS.n1578 394
R1534 VSS.n1583 VSS.n1582 394
R1535 VSS.n1587 VSS.n1586 394
R1536 VSS.n1591 VSS.n1590 394
R1537 VSS.n1595 VSS.n1594 394
R1538 VSS.n1599 VSS.n1598 394
R1539 VSS.n1603 VSS.n1602 394
R1540 VSS.n1607 VSS.n1606 394
R1541 VSS.n1611 VSS.n1610 394
R1542 VSS.n1615 VSS.n1614 394
R1543 VSS.n1619 VSS.n1618 394
R1544 VSS.n1623 VSS.n1622 394
R1545 VSS.n1627 VSS.n1626 394
R1546 VSS.n1631 VSS.n1630 394
R1547 VSS.n1635 VSS.n1634 394
R1548 VSS.n1639 VSS.n1638 394
R1549 VSS.n1643 VSS.n1642 394
R1550 VSS.n1647 VSS.n1646 394
R1551 VSS.n1649 VSS.n1472 394
R1552 VSS.n1653 VSS.n1436 394
R1553 VSS.n1734 VSS.n1433 394
R1554 VSS.n1734 VSS.n1434 394
R1555 VSS.n1434 VSS.n1395 394
R1556 VSS.n1833 VSS.n1395 394
R1557 VSS.n1833 VSS.n1396 394
R1558 VSS.n1407 VSS.n1396 394
R1559 VSS.n1823 VSS.n1407 394
R1560 VSS.n1823 VSS.n1815 394
R1561 VSS.n1815 VSS.n675 394
R1562 VSS.n2169 VSS.n675 394
R1563 VSS.n2169 VSS.n676 394
R1564 VSS.n2165 VSS.n676 394
R1565 VSS.n2165 VSS.n679 394
R1566 VSS.n1327 VSS.n679 394
R1567 VSS.n1330 VSS.n1327 394
R1568 VSS.n1330 VSS.n1324 394
R1569 VSS.n1903 VSS.n1324 394
R1570 VSS.n1903 VSS.n752 394
R1571 VSS.n2148 VSS.n752 394
R1572 VSS.n2148 VSS.n753 394
R1573 VSS.n2144 VSS.n753 394
R1574 VSS.n2144 VSS.n757 394
R1575 VSS.n768 VSS.n757 394
R1576 VSS.n2134 VSS.n768 394
R1577 VSS.n2134 VSS.n769 394
R1578 VSS.n2130 VSS.n769 394
R1579 VSS.n2130 VSS.n772 394
R1580 VSS.n862 VSS.n772 394
R1581 VSS.n2119 VSS.n862 394
R1582 VSS.n2119 VSS.n863 394
R1583 VSS.n1958 VSS.n863 394
R1584 VSS.n1958 VSS.n869 394
R1585 VSS.n2112 VSS.n869 394
R1586 VSS.n2112 VSS.n870 394
R1587 VSS.n881 VSS.n870 394
R1588 VSS.n2102 VSS.n881 394
R1589 VSS.n2102 VSS.n882 394
R1590 VSS.n2096 VSS.n882 394
R1591 VSS.n951 VSS.n950 394
R1592 VSS.n1166 VSS.n950 394
R1593 VSS.n1164 VSS.n1163 394
R1594 VSS.n1160 VSS.n1159 394
R1595 VSS.n1156 VSS.n1155 394
R1596 VSS.n1152 VSS.n1151 394
R1597 VSS.n1148 VSS.n1147 394
R1598 VSS.n1144 VSS.n1143 394
R1599 VSS.n1140 VSS.n1139 394
R1600 VSS.n1136 VSS.n949 394
R1601 VSS.n1133 VSS.n949 394
R1602 VSS.n1131 VSS.n1130 394
R1603 VSS.n1126 VSS.n1124 394
R1604 VSS.n1122 VSS.n956 394
R1605 VSS.n1118 VSS.n1116 394
R1606 VSS.n1114 VSS.n958 394
R1607 VSS.n1110 VSS.n1108 394
R1608 VSS.n1106 VSS.n960 394
R1609 VSS.n1102 VSS.n1100 394
R1610 VSS.n1098 VSS.n962 394
R1611 VSS.n1094 VSS.n1092 394
R1612 VSS.n1090 VSS.n964 394
R1613 VSS.n1086 VSS.n1084 394
R1614 VSS.n1078 VSS.n1076 394
R1615 VSS.n1074 VSS.n968 394
R1616 VSS.n1070 VSS.n1068 394
R1617 VSS.n1066 VSS.n970 394
R1618 VSS.n1062 VSS.n1060 394
R1619 VSS.n1058 VSS.n972 394
R1620 VSS.n1054 VSS.n1052 394
R1621 VSS.n1050 VSS.n974 394
R1622 VSS.n1046 VSS.n1044 394
R1623 VSS.n1042 VSS.n976 394
R1624 VSS.n1038 VSS.n1036 394
R1625 VSS.n1030 VSS.n1028 394
R1626 VSS.n1026 VSS.n980 394
R1627 VSS.n1022 VSS.n1020 394
R1628 VSS.n1018 VSS.n982 394
R1629 VSS.n1014 VSS.n1012 394
R1630 VSS.n1010 VSS.n984 394
R1631 VSS.n1006 VSS.n1004 394
R1632 VSS.n1002 VSS.n986 394
R1633 VSS.n998 VSS.n996 394
R1634 VSS.n994 VSS.n988 394
R1635 VSS.n990 VSS.n887 394
R1636 VSS.n551 VSS.n546 394
R1637 VSS.n555 VSS.n553 394
R1638 VSS.n561 VSS.n544 394
R1639 VSS.n565 VSS.n544 394
R1640 VSS.n565 VSS.n538 394
R1641 VSS.n574 VSS.n538 394
R1642 VSS.n574 VSS.n536 394
R1643 VSS.n578 VSS.n536 394
R1644 VSS.n578 VSS.n446 394
R1645 VSS.n2292 VSS.n446 394
R1646 VSS.n2292 VSS.n447 394
R1647 VSS.n2288 VSS.n447 394
R1648 VSS.n2288 VSS.n450 394
R1649 VSS.n2284 VSS.n450 394
R1650 VSS.n2284 VSS.n455 394
R1651 VSS.n2280 VSS.n455 394
R1652 VSS.n2280 VSS.n457 394
R1653 VSS.n2276 VSS.n457 394
R1654 VSS.n2276 VSS.n462 394
R1655 VSS.n2272 VSS.n462 394
R1656 VSS.n2272 VSS.n464 394
R1657 VSS.n2268 VSS.n464 394
R1658 VSS.n2268 VSS.n469 394
R1659 VSS.n2264 VSS.n469 394
R1660 VSS.n2264 VSS.n471 394
R1661 VSS.n2260 VSS.n471 394
R1662 VSS.n2260 VSS.n476 394
R1663 VSS.n2256 VSS.n476 394
R1664 VSS.n2256 VSS.n478 394
R1665 VSS.n2252 VSS.n478 394
R1666 VSS.n2252 VSS.n483 394
R1667 VSS.n2248 VSS.n483 394
R1668 VSS.n2248 VSS.n485 394
R1669 VSS.n2244 VSS.n485 394
R1670 VSS.n2244 VSS.n490 394
R1671 VSS.n2240 VSS.n490 394
R1672 VSS.n2240 VSS.n492 394
R1673 VSS.n2236 VSS.n492 394
R1674 VSS.n2236 VSS.n497 394
R1675 VSS.n2232 VSS.n497 394
R1676 VSS.n2232 VSS.n499 394
R1677 VSS.n2228 VSS.n499 394
R1678 VSS.n2228 VSS.n504 394
R1679 VSS.n2224 VSS.n504 394
R1680 VSS.n2224 VSS.n506 394
R1681 VSS.n2220 VSS.n506 394
R1682 VSS.n2220 VSS.n511 394
R1683 VSS.n2216 VSS.n511 394
R1684 VSS.n2216 VSS.n513 394
R1685 VSS.n2212 VSS.n513 394
R1686 VSS.n2212 VSS.n518 394
R1687 VSS.n2208 VSS.n518 394
R1688 VSS.n2208 VSS.n520 394
R1689 VSS.n2204 VSS.n520 394
R1690 VSS.n2204 VSS.n525 394
R1691 VSS.n2196 VSS.n529 394
R1692 VSS.n530 VSS.n529 394
R1693 VSS.n559 VSS.n542 394
R1694 VSS.n567 VSS.n542 394
R1695 VSS.n567 VSS.n540 394
R1696 VSS.n572 VSS.n540 394
R1697 VSS.n572 VSS.n534 394
R1698 VSS.n580 VSS.n534 394
R1699 VSS.n581 VSS.n580 394
R1700 VSS.n581 VSS.n444 394
R1701 VSS.n584 VSS.n444 394
R1702 VSS.n584 VSS.n451 394
R1703 VSS.n452 VSS.n451 394
R1704 VSS.n453 VSS.n452 394
R1705 VSS.n589 VSS.n453 394
R1706 VSS.n589 VSS.n458 394
R1707 VSS.n459 VSS.n458 394
R1708 VSS.n460 VSS.n459 394
R1709 VSS.n594 VSS.n460 394
R1710 VSS.n594 VSS.n465 394
R1711 VSS.n466 VSS.n465 394
R1712 VSS.n467 VSS.n466 394
R1713 VSS.n599 VSS.n467 394
R1714 VSS.n599 VSS.n472 394
R1715 VSS.n473 VSS.n472 394
R1716 VSS.n474 VSS.n473 394
R1717 VSS.n604 VSS.n474 394
R1718 VSS.n604 VSS.n479 394
R1719 VSS.n607 VSS.n479 394
R1720 VSS.n607 VSS.n481 394
R1721 VSS.n610 VSS.n481 394
R1722 VSS.n610 VSS.n486 394
R1723 VSS.n487 VSS.n486 394
R1724 VSS.n488 VSS.n487 394
R1725 VSS.n615 VSS.n488 394
R1726 VSS.n615 VSS.n493 394
R1727 VSS.n494 VSS.n493 394
R1728 VSS.n495 VSS.n494 394
R1729 VSS.n620 VSS.n495 394
R1730 VSS.n620 VSS.n500 394
R1731 VSS.n501 VSS.n500 394
R1732 VSS.n502 VSS.n501 394
R1733 VSS.n625 VSS.n502 394
R1734 VSS.n625 VSS.n507 394
R1735 VSS.n508 VSS.n507 394
R1736 VSS.n509 VSS.n508 394
R1737 VSS.n630 VSS.n509 394
R1738 VSS.n630 VSS.n514 394
R1739 VSS.n515 VSS.n514 394
R1740 VSS.n516 VSS.n515 394
R1741 VSS.n635 VSS.n516 394
R1742 VSS.n635 VSS.n521 394
R1743 VSS.n522 VSS.n521 394
R1744 VSS.n523 VSS.n522 394
R1745 VSS.n531 VSS.n523 394
R1746 VSS.n2155 VSS.n702 394
R1747 VSS.n2155 VSS.n703 394
R1748 VSS.n2151 VSS.n703 394
R1749 VSS.n2151 VSS.n748 394
R1750 VSS.n760 VSS.n748 394
R1751 VSS.n2141 VSS.n760 394
R1752 VSS.n2141 VSS.n761 394
R1753 VSS.n2137 VSS.n761 394
R1754 VSS.n2137 VSS.n764 394
R1755 VSS.n776 VSS.n764 394
R1756 VSS.n2127 VSS.n776 394
R1757 VSS.n2123 VSS.n780 394
R1758 VSS.n792 VSS.n780 394
R1759 VSS.n796 VSS.n795 394
R1760 VSS.n800 VSS.n799 394
R1761 VSS.n804 VSS.n803 394
R1762 VSS.n808 VSS.n807 394
R1763 VSS.n812 VSS.n811 394
R1764 VSS.n816 VSS.n815 394
R1765 VSS.n820 VSS.n819 394
R1766 VSS.n824 VSS.n823 394
R1767 VSS.n826 VSS.n791 394
R1768 VSS.n2157 VSS.n696 394
R1769 VSS.n2157 VSS.n699 394
R1770 VSS.n750 VSS.n699 394
R1771 VSS.n839 VSS.n750 394
R1772 VSS.n842 VSS.n839 394
R1773 VSS.n842 VSS.n758 394
R1774 VSS.n830 VSS.n758 394
R1775 VSS.n830 VSS.n766 394
R1776 VSS.n852 VSS.n766 394
R1777 VSS.n853 VSS.n852 394
R1778 VSS.n853 VSS.n774 394
R1779 VSS.n742 VSS.n741 394
R1780 VSS.n738 VSS.n737 394
R1781 VSS.n734 VSS.n733 394
R1782 VSS.n730 VSS.n729 394
R1783 VSS.n726 VSS.n725 394
R1784 VSS.n722 VSS.n721 394
R1785 VSS.n718 VSS.n717 394
R1786 VSS.n714 VSS.n713 394
R1787 VSS.n710 VSS.n709 394
R1788 VSS.n706 VSS.n705 394
R1789 VSS.n2161 VSS.n695 394
R1790 VSS.n2253 VSS.n482 328.791
R1791 VSS.n2247 VSS.n482 328.791
R1792 VSS.n2247 VSS.n2246 328.791
R1793 VSS.n2246 VSS.n2245 328.791
R1794 VSS.n2245 VSS.n489 328.791
R1795 VSS.n2239 VSS.n489 328.791
R1796 VSS.n2239 VSS.n2238 328.791
R1797 VSS.n2238 VSS.n2237 328.791
R1798 VSS.n2237 VSS.n496 328.791
R1799 VSS.n2231 VSS.n496 328.791
R1800 VSS.n2231 VSS.n2230 328.791
R1801 VSS.n2230 VSS.n2229 328.791
R1802 VSS.n2229 VSS.n503 328.791
R1803 VSS.n2223 VSS.n503 328.791
R1804 VSS.n2223 VSS.n2222 328.791
R1805 VSS.n2222 VSS.n2221 328.791
R1806 VSS.n2221 VSS.n510 328.791
R1807 VSS.n2215 VSS.n510 328.791
R1808 VSS.n2215 VSS.n2214 328.791
R1809 VSS.n2214 VSS.n2213 328.791
R1810 VSS.n2213 VSS.n517 328.791
R1811 VSS.n2207 VSS.n517 328.791
R1812 VSS.n2207 VSS.n2206 328.791
R1813 VSS.n2206 VSS.n2205 328.791
R1814 VSS.n2205 VSS.n524 328.791
R1815 VSS.n71 VSS.n70 325.69
R1816 VSS.n16 VSS.n11 325.69
R1817 VSS.n1518 VSS.n1438 269.089
R1818 VSS.n1515 VSS.n1438 269.089
R1819 VSS.n2556 VSS.n98 261
R1820 VSS.n932 VSS.t103 259.252
R1821 VSS.n1292 VSS.t62 259.252
R1822 VSS.n1837 VSS.t69 259.252
R1823 VSS.n1883 VSS.t66 259.252
R1824 VSS.n1236 VSS.t106 258.99
R1825 VSS.n1237 VSS.t91 258.99
R1826 VSS.n1238 VSS.t75 258.99
R1827 VSS.n1239 VSS.t123 258.99
R1828 VSS.n1242 VSS.t111 258.99
R1829 VSS.n1241 VSS.t115 258.99
R1830 VSS.n1240 VSS.t97 258.99
R1831 VSS.n1195 VSS.t77 258.99
R1832 VSS.n1374 VSS.t101 258.99
R1833 VSS.n1387 VSS.t125 258.99
R1834 VSS.n1388 VSS.t60 258.99
R1835 VSS.n1389 VSS.t64 258.99
R1836 VSS.n1882 VSS.t113 258.99
R1837 VSS.n1881 VSS.t93 258.99
R1838 VSS.n1880 VSS.t95 258.99
R1839 VSS.n1879 VSS.t99 258.99
R1840 VSS.n1276 VSS.n1246 253.042
R1841 VSS.n1209 VSS.n1208 253.042
R1842 VSS.n1371 VSS.n1370 253.042
R1843 VSS.n1849 VSS.n1847 253.042
R1844 VSS.n554 VSS.n547 218.815
R1845 VSS.n552 VSS.n547 218.815
R1846 VSS.n2195 VSS.n2193 218.815
R1847 VSS.n2193 VSS.n643 218.815
R1848 VSS.n1173 VSS.n1172 218.815
R1849 VSS.n1173 VSS.n941 218.815
R1850 VSS.n1173 VSS.n942 218.815
R1851 VSS.n1173 VSS.n943 218.815
R1852 VSS.n1173 VSS.n944 218.815
R1853 VSS.n1173 VSS.n945 218.815
R1854 VSS.n1173 VSS.n946 218.815
R1855 VSS.n1173 VSS.n947 218.815
R1856 VSS.n1173 VSS.n948 218.815
R1857 VSS.n2192 VSS.n653 218.815
R1858 VSS.n2192 VSS.n652 218.815
R1859 VSS.n2192 VSS.n651 218.815
R1860 VSS.n2192 VSS.n650 218.815
R1861 VSS.n2192 VSS.n649 218.815
R1862 VSS.n2192 VSS.n648 218.815
R1863 VSS.n2192 VSS.n647 218.815
R1864 VSS.n2192 VSS.n646 218.815
R1865 VSS.n2192 VSS.n645 218.815
R1866 VSS.n2192 VSS.n644 218.815
R1867 VSS.n1807 VSS.n680 218.815
R1868 VSS.n1800 VSS.n680 218.815
R1869 VSS.n1798 VSS.n680 218.815
R1870 VSS.n1792 VSS.n680 218.815
R1871 VSS.n1790 VSS.n680 218.815
R1872 VSS.n1784 VSS.n680 218.815
R1873 VSS.n1782 VSS.n680 218.815
R1874 VSS.n1776 VSS.n680 218.815
R1875 VSS.n1774 VSS.n680 218.815
R1876 VSS.n1768 VSS.n680 218.815
R1877 VSS.n1766 VSS.n680 218.815
R1878 VSS.n1680 VSS.n98 218.815
R1879 VSS.n1686 VSS.n98 218.815
R1880 VSS.n1672 VSS.n98 218.815
R1881 VSS.n1693 VSS.n98 218.815
R1882 VSS.n1669 VSS.n98 218.815
R1883 VSS.n1700 VSS.n98 218.815
R1884 VSS.n1666 VSS.n98 218.815
R1885 VSS.n1707 VSS.n98 218.815
R1886 VSS.n1663 VSS.n98 218.815
R1887 VSS.n1714 VSS.n98 218.815
R1888 VSS.n1717 VSS.n98 218.815
R1889 VSS.n2080 VSS.n2079 218.815
R1890 VSS.n2079 VSS.n903 218.815
R1891 VSS.n2079 VSS.n904 218.815
R1892 VSS.n2079 VSS.n905 218.815
R1893 VSS.n2079 VSS.n906 218.815
R1894 VSS.n2079 VSS.n907 218.815
R1895 VSS.n2079 VSS.n908 218.815
R1896 VSS.n2079 VSS.n909 218.815
R1897 VSS.n2079 VSS.n910 218.815
R1898 VSS.n2079 VSS.n911 218.815
R1899 VSS.n2079 VSS.n912 218.815
R1900 VSS.n2014 VSS.n2013 218.815
R1901 VSS.n2013 VSS.n1960 218.815
R1902 VSS.n2013 VSS.n1961 218.815
R1903 VSS.n2013 VSS.n1962 218.815
R1904 VSS.n2013 VSS.n1963 218.815
R1905 VSS.n2013 VSS.n1964 218.815
R1906 VSS.n2013 VSS.n1965 218.815
R1907 VSS.n2013 VSS.n1966 218.815
R1908 VSS.n2013 VSS.n1967 218.815
R1909 VSS.n2013 VSS.n1968 218.815
R1910 VSS.n2013 VSS.n1969 218.815
R1911 VSS.n2556 VSS.n2555 218.815
R1912 VSS.n2556 VSS.n81 218.815
R1913 VSS.n2556 VSS.n82 218.815
R1914 VSS.n2556 VSS.n83 218.815
R1915 VSS.n2556 VSS.n84 218.815
R1916 VSS.n2556 VSS.n85 218.815
R1917 VSS.n2556 VSS.n86 218.815
R1918 VSS.n2556 VSS.n87 218.815
R1919 VSS.n2556 VSS.n88 218.815
R1920 VSS.n2556 VSS.n89 218.815
R1921 VSS.n2556 VSS.n90 218.815
R1922 VSS.n2557 VSS.n2556 218.815
R1923 VSS.n2556 VSS.n91 218.815
R1924 VSS.n2556 VSS.n92 218.815
R1925 VSS.n2556 VSS.n93 218.815
R1926 VSS.n2556 VSS.n94 218.815
R1927 VSS.n2556 VSS.n95 218.815
R1928 VSS.n2556 VSS.n96 218.815
R1929 VSS.n2556 VSS.n97 218.815
R1930 VSS.n425 VSS.n220 218.815
R1931 VSS.n423 VSS.n220 218.815
R1932 VSS.n417 VSS.n220 218.815
R1933 VSS.n415 VSS.n220 218.815
R1934 VSS.n409 VSS.n220 218.815
R1935 VSS.n407 VSS.n220 218.815
R1936 VSS.n401 VSS.n220 218.815
R1937 VSS.n399 VSS.n220 218.815
R1938 VSS.n290 VSS.n220 218.815
R1939 VSS.n288 VSS.n220 218.815
R1940 VSS.n278 VSS.n220 218.815
R1941 VSS.n276 VSS.n220 218.815
R1942 VSS.n268 VSS.n220 218.815
R1943 VSS.n266 VSS.n220 218.815
R1944 VSS.n260 VSS.n220 218.815
R1945 VSS.n258 VSS.n220 218.815
R1946 VSS.n252 VSS.n220 218.815
R1947 VSS.n250 VSS.n220 218.815
R1948 VSS.n244 VSS.n220 218.815
R1949 VSS.n1132 VSS.n890 218.815
R1950 VSS.n1125 VSS.n890 218.815
R1951 VSS.n1123 VSS.n890 218.815
R1952 VSS.n1117 VSS.n890 218.815
R1953 VSS.n1115 VSS.n890 218.815
R1954 VSS.n1109 VSS.n890 218.815
R1955 VSS.n1107 VSS.n890 218.815
R1956 VSS.n1101 VSS.n890 218.815
R1957 VSS.n1099 VSS.n890 218.815
R1958 VSS.n1093 VSS.n890 218.815
R1959 VSS.n1091 VSS.n890 218.815
R1960 VSS.n1085 VSS.n890 218.815
R1961 VSS.n1083 VSS.n890 218.815
R1962 VSS.n1077 VSS.n890 218.815
R1963 VSS.n1075 VSS.n890 218.815
R1964 VSS.n1069 VSS.n890 218.815
R1965 VSS.n1067 VSS.n890 218.815
R1966 VSS.n1061 VSS.n890 218.815
R1967 VSS.n1059 VSS.n890 218.815
R1968 VSS.n1053 VSS.n890 218.815
R1969 VSS.n1051 VSS.n890 218.815
R1970 VSS.n1045 VSS.n890 218.815
R1971 VSS.n1043 VSS.n890 218.815
R1972 VSS.n1037 VSS.n890 218.815
R1973 VSS.n1035 VSS.n890 218.815
R1974 VSS.n1029 VSS.n890 218.815
R1975 VSS.n1027 VSS.n890 218.815
R1976 VSS.n1021 VSS.n890 218.815
R1977 VSS.n1019 VSS.n890 218.815
R1978 VSS.n1013 VSS.n890 218.815
R1979 VSS.n1011 VSS.n890 218.815
R1980 VSS.n1005 VSS.n890 218.815
R1981 VSS.n1003 VSS.n890 218.815
R1982 VSS.n997 VSS.n890 218.815
R1983 VSS.n995 VSS.n890 218.815
R1984 VSS.n989 VSS.n890 218.815
R1985 VSS.n1725 VSS.n1724 218.815
R1986 VSS.n1724 VSS.n1654 218.815
R1987 VSS.n1724 VSS.n1471 218.815
R1988 VSS.n1724 VSS.n1470 218.815
R1989 VSS.n1724 VSS.n1469 218.815
R1990 VSS.n1724 VSS.n1468 218.815
R1991 VSS.n1724 VSS.n1467 218.815
R1992 VSS.n1724 VSS.n1466 218.815
R1993 VSS.n1724 VSS.n1465 218.815
R1994 VSS.n1724 VSS.n1464 218.815
R1995 VSS.n1724 VSS.n1463 218.815
R1996 VSS.n1724 VSS.n1461 218.815
R1997 VSS.n1724 VSS.n1460 218.815
R1998 VSS.n1724 VSS.n1459 218.815
R1999 VSS.n1724 VSS.n1458 218.815
R2000 VSS.n1724 VSS.n1457 218.815
R2001 VSS.n1724 VSS.n1456 218.815
R2002 VSS.n1724 VSS.n1455 218.815
R2003 VSS.n1724 VSS.n1454 218.815
R2004 VSS.n1724 VSS.n1453 218.815
R2005 VSS.n1724 VSS.n1452 218.815
R2006 VSS.n1724 VSS.n1451 218.815
R2007 VSS.n1724 VSS.n1449 218.815
R2008 VSS.n1724 VSS.n1448 218.815
R2009 VSS.n1724 VSS.n1447 218.815
R2010 VSS.n1724 VSS.n1446 218.815
R2011 VSS.n1724 VSS.n1445 218.815
R2012 VSS.n1724 VSS.n1444 218.815
R2013 VSS.n1724 VSS.n1443 218.815
R2014 VSS.n1724 VSS.n1442 218.815
R2015 VSS.n1724 VSS.n1441 218.815
R2016 VSS.n1724 VSS.n1440 218.815
R2017 VSS.n1724 VSS.n1439 218.815
R2018 VSS.n1724 VSS.n1437 218.815
R2019 VSS.n2162 VSS.n693 218.815
R2020 VSS.n2162 VSS.n692 218.815
R2021 VSS.n2162 VSS.n691 218.815
R2022 VSS.n2162 VSS.n690 218.815
R2023 VSS.n2162 VSS.n689 218.815
R2024 VSS.n2162 VSS.n688 218.815
R2025 VSS.n2162 VSS.n687 218.815
R2026 VSS.n2162 VSS.n686 218.815
R2027 VSS.n2162 VSS.n685 218.815
R2028 VSS.n2162 VSS.n684 218.815
R2029 VSS.n2162 VSS.n683 218.815
R2030 VSS.n2122 VSS.n2121 218.815
R2031 VSS.n2121 VSS.n782 218.815
R2032 VSS.n2121 VSS.n783 218.815
R2033 VSS.n2121 VSS.n784 218.815
R2034 VSS.n2121 VSS.n785 218.815
R2035 VSS.n2121 VSS.n786 218.815
R2036 VSS.n2121 VSS.n787 218.815
R2037 VSS.n2121 VSS.n788 218.815
R2038 VSS.n2121 VSS.n789 218.815
R2039 VSS.n2121 VSS.n790 218.815
R2040 VSS.n2121 VSS.n858 218.815
R2041 VSS.n1566 VSS.n1450 198.87
R2042 VSS.n1614 VSS.n1462 198.87
R2043 VSS.n1611 VSS.n1462 198.87
R2044 VSS.n1563 VSS.n1450 198.87
R2045 VSS.n1724 VSS.n1462 193.066
R2046 VSS.n1724 VSS.n1450 193.066
R2047 VSS.n560 VSS.n547 185.895
R2048 VSS.n328 VSS.n327 185
R2049 VSS.n328 VSS.n300 185
R2050 VSS.n330 VSS.n329 185
R2051 VSS.n329 VSS.n298 185
R2052 VSS.n312 VSS.n304 185
R2053 VSS.n312 VSS.n303 185
R2054 VSS.n313 VSS.n312 185
R2055 VSS.n390 VSS.n389 185
R2056 VSS.n389 VSS.n373 185
R2057 VSS.n388 VSS.n387 185
R2058 VSS.n388 VSS.n375 185
R2059 VSS.n367 VSS.n359 185
R2060 VSS.n367 VSS.n358 185
R2061 VSS.n368 VSS.n367 185
R2062 VSS.n70 VSS.n69 185
R2063 VSS.n47 VSS.n46 185
R2064 VSS.n64 VSS.n63 185
R2065 VSS.n58 VSS.n57 185
R2066 VSS.n58 VSS.n50 185
R2067 VSS.n30 VSS.n29 185
R2068 VSS.n29 VSS.n28 185
R2069 VSS.n16 VSS.n15 185
R2070 VSS.n18 VSS.n17 185
R2071 VSS.n20 VSS.n8 185
R2072 VSS.n1277 VSS.n1276 185
R2073 VSS.n1275 VSS.n1274 185
R2074 VSS.n1250 VSS.n1249 185
R2075 VSS.n1269 VSS.n1268 185
R2076 VSS.n1267 VSS.n1266 185
R2077 VSS.n1254 VSS.n1253 185
R2078 VSS.n1261 VSS.n1260 185
R2079 VSS.n1259 VSS.n1258 185
R2080 VSS.n1210 VSS.n1209 185
R2081 VSS.n1205 VSS.n1204 185
R2082 VSS.n1216 VSS.n1215 185
R2083 VSS.n1218 VSS.n1217 185
R2084 VSS.n1201 VSS.n1200 185
R2085 VSS.n1225 VSS.n1224 185
R2086 VSS.n1227 VSS.n1226 185
R2087 VSS.n1229 VSS.n1197 185
R2088 VSS.n1349 VSS.n1348 185
R2089 VSS.n1354 VSS.n1353 185
R2090 VSS.n1356 VSS.n1355 185
R2091 VSS.n1345 VSS.n1344 185
R2092 VSS.n1362 VSS.n1361 185
R2093 VSS.n1364 VSS.n1363 185
R2094 VSS.n1341 VSS.n1340 185
R2095 VSS.n1370 VSS.n1369 185
R2096 VSS.n1871 VSS.n1870 185
R2097 VSS.n1840 VSS.n1839 185
R2098 VSS.n1865 VSS.n1864 185
R2099 VSS.n1863 VSS.n1862 185
R2100 VSS.n1844 VSS.n1843 185
R2101 VSS.n1857 VSS.n1856 185
R2102 VSS.n1855 VSS.n1854 185
R2103 VSS.n1848 VSS.n1847 185
R2104 VSS.n1257 VSS.t105 178.418
R2105 VSS.t63 VSS.n1230 178.418
R2106 VSS.n1350 VSS.t68 178.418
R2107 VSS.t70 VSS.n1838 178.418
R2108 VSS.t110 VSS.n62 175.332
R2109 VSS.t120 VSS.n21 175.332
R2110 VSS.n2192 VSS.n2191 163.94
R2111 VSS.n1174 VSS.n1173 163.94
R2112 VSS.n1724 VSS.n1438 157.957
R2113 VSS.n244 VSS.n243 147.374
R2114 VSS.n251 VSS.n250 147.374
R2115 VSS.n252 VSS.n241 147.374
R2116 VSS.n259 VSS.n258 147.374
R2117 VSS.n260 VSS.n239 147.374
R2118 VSS.n267 VSS.n266 147.374
R2119 VSS.n268 VSS.n237 147.374
R2120 VSS.n277 VSS.n276 147.374
R2121 VSS.n278 VSS.n233 147.374
R2122 VSS.n289 VSS.n288 147.374
R2123 VSS.n290 VSS.n229 147.374
R2124 VSS.n400 VSS.n399 147.374
R2125 VSS.n401 VSS.n227 147.374
R2126 VSS.n408 VSS.n407 147.374
R2127 VSS.n409 VSS.n225 147.374
R2128 VSS.n416 VSS.n415 147.374
R2129 VSS.n417 VSS.n223 147.374
R2130 VSS.n424 VSS.n423 147.374
R2131 VSS.n425 VSS.n221 147.374
R2132 VSS.n2555 VSS.n2554 147.374
R2133 VSS.n2549 VSS.n81 147.374
R2134 VSS.n2546 VSS.n82 147.374
R2135 VSS.n2542 VSS.n83 147.374
R2136 VSS.n2538 VSS.n84 147.374
R2137 VSS.n2534 VSS.n85 147.374
R2138 VSS.n2530 VSS.n86 147.374
R2139 VSS.n2526 VSS.n87 147.374
R2140 VSS.n2519 VSS.n88 147.374
R2141 VSS.n2515 VSS.n89 147.374
R2142 VSS.n2505 VSS.n90 147.374
R2143 VSS.n2557 VSS.n79 147.374
R2144 VSS.n91 VSS.n78 147.374
R2145 VSS.n2468 VSS.n92 147.374
R2146 VSS.n2472 VSS.n93 147.374
R2147 VSS.n2476 VSS.n94 147.374
R2148 VSS.n2480 VSS.n95 147.374
R2149 VSS.n2484 VSS.n96 147.374
R2150 VSS.n2488 VSS.n97 147.374
R2151 VSS.n2008 VSS.n1969 147.374
R2152 VSS.n2004 VSS.n1968 147.374
R2153 VSS.n2000 VSS.n1967 147.374
R2154 VSS.n1996 VSS.n1966 147.374
R2155 VSS.n1992 VSS.n1965 147.374
R2156 VSS.n1988 VSS.n1964 147.374
R2157 VSS.n1984 VSS.n1963 147.374
R2158 VSS.n1980 VSS.n1962 147.374
R2159 VSS.n1976 VSS.n1961 147.374
R2160 VSS.n1972 VSS.n1960 147.374
R2161 VSS.n2015 VSS.n2014 147.374
R2162 VSS.n2081 VSS.n2080 147.374
R2163 VSS.n913 VSS.n903 147.374
R2164 VSS.n2073 VSS.n904 147.374
R2165 VSS.n2069 VSS.n905 147.374
R2166 VSS.n919 VSS.n906 147.374
R2167 VSS.n2061 VSS.n907 147.374
R2168 VSS.n2057 VSS.n908 147.374
R2169 VSS.n2052 VSS.n909 147.374
R2170 VSS.n2048 VSS.n910 147.374
R2171 VSS.n2044 VSS.n911 147.374
R2172 VSS.n2040 VSS.n912 147.374
R2173 VSS.n1717 VSS.n1716 147.374
R2174 VSS.n1714 VSS.n1713 147.374
R2175 VSS.n1709 VSS.n1663 147.374
R2176 VSS.n1707 VSS.n1706 147.374
R2177 VSS.n1702 VSS.n1666 147.374
R2178 VSS.n1700 VSS.n1699 147.374
R2179 VSS.n1695 VSS.n1669 147.374
R2180 VSS.n1693 VSS.n1692 147.374
R2181 VSS.n1688 VSS.n1672 147.374
R2182 VSS.n1686 VSS.n1685 147.374
R2183 VSS.n1681 VSS.n1680 147.374
R2184 VSS.n1808 VSS.n1807 147.374
R2185 VSS.n1800 VSS.n1412 147.374
R2186 VSS.n1799 VSS.n1798 147.374
R2187 VSS.n1792 VSS.n1414 147.374
R2188 VSS.n1791 VSS.n1790 147.374
R2189 VSS.n1784 VSS.n1416 147.374
R2190 VSS.n1783 VSS.n1782 147.374
R2191 VSS.n1776 VSS.n1418 147.374
R2192 VSS.n1775 VSS.n1774 147.374
R2193 VSS.n1768 VSS.n1420 147.374
R2194 VSS.n1767 VSS.n1766 147.374
R2195 VSS.n1474 VSS.n644 147.374
R2196 VSS.n1478 VSS.n645 147.374
R2197 VSS.n1482 VSS.n646 147.374
R2198 VSS.n1486 VSS.n647 147.374
R2199 VSS.n1490 VSS.n648 147.374
R2200 VSS.n1494 VSS.n649 147.374
R2201 VSS.n1498 VSS.n650 147.374
R2202 VSS.n1502 VSS.n651 147.374
R2203 VSS.n1506 VSS.n652 147.374
R2204 VSS.n1510 VSS.n653 147.374
R2205 VSS.n1514 VSS.n1437 147.374
R2206 VSS.n1522 VSS.n1439 147.374
R2207 VSS.n1526 VSS.n1440 147.374
R2208 VSS.n1530 VSS.n1441 147.374
R2209 VSS.n1534 VSS.n1442 147.374
R2210 VSS.n1538 VSS.n1443 147.374
R2211 VSS.n1542 VSS.n1444 147.374
R2212 VSS.n1546 VSS.n1445 147.374
R2213 VSS.n1550 VSS.n1446 147.374
R2214 VSS.n1554 VSS.n1447 147.374
R2215 VSS.n1558 VSS.n1448 147.374
R2216 VSS.n1562 VSS.n1449 147.374
R2217 VSS.n1570 VSS.n1451 147.374
R2218 VSS.n1574 VSS.n1452 147.374
R2219 VSS.n1578 VSS.n1453 147.374
R2220 VSS.n1582 VSS.n1454 147.374
R2221 VSS.n1586 VSS.n1455 147.374
R2222 VSS.n1590 VSS.n1456 147.374
R2223 VSS.n1594 VSS.n1457 147.374
R2224 VSS.n1598 VSS.n1458 147.374
R2225 VSS.n1602 VSS.n1459 147.374
R2226 VSS.n1606 VSS.n1460 147.374
R2227 VSS.n1610 VSS.n1461 147.374
R2228 VSS.n1618 VSS.n1463 147.374
R2229 VSS.n1622 VSS.n1464 147.374
R2230 VSS.n1626 VSS.n1465 147.374
R2231 VSS.n1630 VSS.n1466 147.374
R2232 VSS.n1634 VSS.n1467 147.374
R2233 VSS.n1638 VSS.n1468 147.374
R2234 VSS.n1642 VSS.n1469 147.374
R2235 VSS.n1646 VSS.n1470 147.374
R2236 VSS.n1649 VSS.n1471 147.374
R2237 VSS.n1654 VSS.n1653 147.374
R2238 VSS.n1726 VSS.n1725 147.374
R2239 VSS.n1172 VSS.n1171 147.374
R2240 VSS.n1166 VSS.n941 147.374
R2241 VSS.n1163 VSS.n942 147.374
R2242 VSS.n1159 VSS.n943 147.374
R2243 VSS.n1155 VSS.n944 147.374
R2244 VSS.n1151 VSS.n945 147.374
R2245 VSS.n1147 VSS.n946 147.374
R2246 VSS.n1143 VSS.n947 147.374
R2247 VSS.n1139 VSS.n948 147.374
R2248 VSS.n1133 VSS.n1132 147.374
R2249 VSS.n1125 VSS.n954 147.374
R2250 VSS.n1124 VSS.n1123 147.374
R2251 VSS.n1117 VSS.n956 147.374
R2252 VSS.n1116 VSS.n1115 147.374
R2253 VSS.n1109 VSS.n958 147.374
R2254 VSS.n1108 VSS.n1107 147.374
R2255 VSS.n1101 VSS.n960 147.374
R2256 VSS.n1100 VSS.n1099 147.374
R2257 VSS.n1093 VSS.n962 147.374
R2258 VSS.n1092 VSS.n1091 147.374
R2259 VSS.n1085 VSS.n964 147.374
R2260 VSS.n1084 VSS.n1083 147.374
R2261 VSS.n1077 VSS.n966 147.374
R2262 VSS.n1076 VSS.n1075 147.374
R2263 VSS.n1069 VSS.n968 147.374
R2264 VSS.n1068 VSS.n1067 147.374
R2265 VSS.n1061 VSS.n970 147.374
R2266 VSS.n1060 VSS.n1059 147.374
R2267 VSS.n1053 VSS.n972 147.374
R2268 VSS.n1052 VSS.n1051 147.374
R2269 VSS.n1045 VSS.n974 147.374
R2270 VSS.n1044 VSS.n1043 147.374
R2271 VSS.n1037 VSS.n976 147.374
R2272 VSS.n1036 VSS.n1035 147.374
R2273 VSS.n1029 VSS.n978 147.374
R2274 VSS.n1028 VSS.n1027 147.374
R2275 VSS.n1021 VSS.n980 147.374
R2276 VSS.n1020 VSS.n1019 147.374
R2277 VSS.n1013 VSS.n982 147.374
R2278 VSS.n1012 VSS.n1011 147.374
R2279 VSS.n1005 VSS.n984 147.374
R2280 VSS.n1004 VSS.n1003 147.374
R2281 VSS.n997 VSS.n986 147.374
R2282 VSS.n996 VSS.n995 147.374
R2283 VSS.n989 VSS.n988 147.374
R2284 VSS.n553 VSS.n552 147.374
R2285 VSS.n554 VSS.n548 147.374
R2286 VSS.n2195 VSS.n2194 147.374
R2287 VSS.n643 VSS.n530 147.374
R2288 VSS.n555 VSS.n554 147.374
R2289 VSS.n552 VSS.n551 147.374
R2290 VSS.n2196 VSS.n2195 147.374
R2291 VSS.n643 VSS.n642 147.374
R2292 VSS.n1172 VSS.n951 147.374
R2293 VSS.n1164 VSS.n941 147.374
R2294 VSS.n1160 VSS.n942 147.374
R2295 VSS.n1156 VSS.n943 147.374
R2296 VSS.n1152 VSS.n944 147.374
R2297 VSS.n1148 VSS.n945 147.374
R2298 VSS.n1144 VSS.n946 147.374
R2299 VSS.n1140 VSS.n947 147.374
R2300 VSS.n1136 VSS.n948 147.374
R2301 VSS.n1507 VSS.n653 147.374
R2302 VSS.n1503 VSS.n652 147.374
R2303 VSS.n1499 VSS.n651 147.374
R2304 VSS.n1495 VSS.n650 147.374
R2305 VSS.n1491 VSS.n649 147.374
R2306 VSS.n1487 VSS.n648 147.374
R2307 VSS.n1483 VSS.n647 147.374
R2308 VSS.n1479 VSS.n646 147.374
R2309 VSS.n1475 VSS.n645 147.374
R2310 VSS.n655 VSS.n644 147.374
R2311 VSS.n1807 VSS.n1806 147.374
R2312 VSS.n1801 VSS.n1800 147.374
R2313 VSS.n1798 VSS.n1797 147.374
R2314 VSS.n1793 VSS.n1792 147.374
R2315 VSS.n1790 VSS.n1789 147.374
R2316 VSS.n1785 VSS.n1784 147.374
R2317 VSS.n1782 VSS.n1781 147.374
R2318 VSS.n1777 VSS.n1776 147.374
R2319 VSS.n1774 VSS.n1773 147.374
R2320 VSS.n1769 VSS.n1768 147.374
R2321 VSS.n1766 VSS.n1765 147.374
R2322 VSS.n1680 VSS.n1673 147.374
R2323 VSS.n1687 VSS.n1686 147.374
R2324 VSS.n1672 VSS.n1670 147.374
R2325 VSS.n1694 VSS.n1693 147.374
R2326 VSS.n1669 VSS.n1667 147.374
R2327 VSS.n1701 VSS.n1700 147.374
R2328 VSS.n1666 VSS.n1664 147.374
R2329 VSS.n1708 VSS.n1707 147.374
R2330 VSS.n1663 VSS.n1661 147.374
R2331 VSS.n1715 VSS.n1714 147.374
R2332 VSS.n1718 VSS.n1717 147.374
R2333 VSS.n2080 VSS.n902 147.374
R2334 VSS.n2074 VSS.n903 147.374
R2335 VSS.n2070 VSS.n904 147.374
R2336 VSS.n918 VSS.n905 147.374
R2337 VSS.n2062 VSS.n906 147.374
R2338 VSS.n2058 VSS.n907 147.374
R2339 VSS.n2053 VSS.n908 147.374
R2340 VSS.n2049 VSS.n909 147.374
R2341 VSS.n2045 VSS.n910 147.374
R2342 VSS.n2041 VSS.n911 147.374
R2343 VSS.n2037 VSS.n912 147.374
R2344 VSS.n2014 VSS.n925 147.374
R2345 VSS.n1975 VSS.n1960 147.374
R2346 VSS.n1979 VSS.n1961 147.374
R2347 VSS.n1983 VSS.n1962 147.374
R2348 VSS.n1987 VSS.n1963 147.374
R2349 VSS.n1991 VSS.n1964 147.374
R2350 VSS.n1995 VSS.n1965 147.374
R2351 VSS.n1999 VSS.n1966 147.374
R2352 VSS.n2003 VSS.n1967 147.374
R2353 VSS.n2007 VSS.n1968 147.374
R2354 VSS.n1970 VSS.n1969 147.374
R2355 VSS.n2555 VSS.n100 147.374
R2356 VSS.n2547 VSS.n81 147.374
R2357 VSS.n2543 VSS.n82 147.374
R2358 VSS.n2539 VSS.n83 147.374
R2359 VSS.n2535 VSS.n84 147.374
R2360 VSS.n2531 VSS.n85 147.374
R2361 VSS.n2527 VSS.n86 147.374
R2362 VSS.n2518 VSS.n87 147.374
R2363 VSS.n2516 VSS.n88 147.374
R2364 VSS.n2504 VSS.n89 147.374
R2365 VSS.n2508 VSS.n90 147.374
R2366 VSS.n2558 VSS.n2557 147.374
R2367 VSS.n2467 VSS.n91 147.374
R2368 VSS.n2471 VSS.n92 147.374
R2369 VSS.n2475 VSS.n93 147.374
R2370 VSS.n2479 VSS.n94 147.374
R2371 VSS.n2483 VSS.n95 147.374
R2372 VSS.n2487 VSS.n96 147.374
R2373 VSS.n2490 VSS.n97 147.374
R2374 VSS.n426 VSS.n425 147.374
R2375 VSS.n423 VSS.n422 147.374
R2376 VSS.n418 VSS.n417 147.374
R2377 VSS.n415 VSS.n414 147.374
R2378 VSS.n410 VSS.n409 147.374
R2379 VSS.n407 VSS.n406 147.374
R2380 VSS.n402 VSS.n401 147.374
R2381 VSS.n399 VSS.n398 147.374
R2382 VSS.n291 VSS.n290 147.374
R2383 VSS.n288 VSS.n287 147.374
R2384 VSS.n279 VSS.n278 147.374
R2385 VSS.n276 VSS.n275 147.374
R2386 VSS.n269 VSS.n268 147.374
R2387 VSS.n266 VSS.n265 147.374
R2388 VSS.n261 VSS.n260 147.374
R2389 VSS.n258 VSS.n257 147.374
R2390 VSS.n253 VSS.n252 147.374
R2391 VSS.n250 VSS.n249 147.374
R2392 VSS.n245 VSS.n244 147.374
R2393 VSS.n1132 VSS.n1131 147.374
R2394 VSS.n1126 VSS.n1125 147.374
R2395 VSS.n1123 VSS.n1122 147.374
R2396 VSS.n1118 VSS.n1117 147.374
R2397 VSS.n1115 VSS.n1114 147.374
R2398 VSS.n1110 VSS.n1109 147.374
R2399 VSS.n1107 VSS.n1106 147.374
R2400 VSS.n1102 VSS.n1101 147.374
R2401 VSS.n1099 VSS.n1098 147.374
R2402 VSS.n1094 VSS.n1093 147.374
R2403 VSS.n1091 VSS.n1090 147.374
R2404 VSS.n1086 VSS.n1085 147.374
R2405 VSS.n1083 VSS.n1082 147.374
R2406 VSS.n1078 VSS.n1077 147.374
R2407 VSS.n1075 VSS.n1074 147.374
R2408 VSS.n1070 VSS.n1069 147.374
R2409 VSS.n1067 VSS.n1066 147.374
R2410 VSS.n1062 VSS.n1061 147.374
R2411 VSS.n1059 VSS.n1058 147.374
R2412 VSS.n1054 VSS.n1053 147.374
R2413 VSS.n1051 VSS.n1050 147.374
R2414 VSS.n1046 VSS.n1045 147.374
R2415 VSS.n1043 VSS.n1042 147.374
R2416 VSS.n1038 VSS.n1037 147.374
R2417 VSS.n1035 VSS.n1034 147.374
R2418 VSS.n1030 VSS.n1029 147.374
R2419 VSS.n1027 VSS.n1026 147.374
R2420 VSS.n1022 VSS.n1021 147.374
R2421 VSS.n1019 VSS.n1018 147.374
R2422 VSS.n1014 VSS.n1013 147.374
R2423 VSS.n1011 VSS.n1010 147.374
R2424 VSS.n1006 VSS.n1005 147.374
R2425 VSS.n1003 VSS.n1002 147.374
R2426 VSS.n998 VSS.n997 147.374
R2427 VSS.n995 VSS.n994 147.374
R2428 VSS.n990 VSS.n989 147.374
R2429 VSS.n1725 VSS.n1436 147.374
R2430 VSS.n1654 VSS.n1472 147.374
R2431 VSS.n1647 VSS.n1471 147.374
R2432 VSS.n1643 VSS.n1470 147.374
R2433 VSS.n1639 VSS.n1469 147.374
R2434 VSS.n1635 VSS.n1468 147.374
R2435 VSS.n1631 VSS.n1467 147.374
R2436 VSS.n1627 VSS.n1466 147.374
R2437 VSS.n1623 VSS.n1465 147.374
R2438 VSS.n1619 VSS.n1464 147.374
R2439 VSS.n1615 VSS.n1463 147.374
R2440 VSS.n1607 VSS.n1461 147.374
R2441 VSS.n1603 VSS.n1460 147.374
R2442 VSS.n1599 VSS.n1459 147.374
R2443 VSS.n1595 VSS.n1458 147.374
R2444 VSS.n1591 VSS.n1457 147.374
R2445 VSS.n1587 VSS.n1456 147.374
R2446 VSS.n1583 VSS.n1455 147.374
R2447 VSS.n1579 VSS.n1454 147.374
R2448 VSS.n1575 VSS.n1453 147.374
R2449 VSS.n1571 VSS.n1452 147.374
R2450 VSS.n1567 VSS.n1451 147.374
R2451 VSS.n1559 VSS.n1449 147.374
R2452 VSS.n1555 VSS.n1448 147.374
R2453 VSS.n1551 VSS.n1447 147.374
R2454 VSS.n1547 VSS.n1446 147.374
R2455 VSS.n1543 VSS.n1445 147.374
R2456 VSS.n1539 VSS.n1444 147.374
R2457 VSS.n1535 VSS.n1443 147.374
R2458 VSS.n1531 VSS.n1442 147.374
R2459 VSS.n1527 VSS.n1441 147.374
R2460 VSS.n1523 VSS.n1440 147.374
R2461 VSS.n1519 VSS.n1439 147.374
R2462 VSS.n1511 VSS.n1437 147.374
R2463 VSS.n2122 VSS.n777 147.374
R2464 VSS.n792 VSS.n782 147.374
R2465 VSS.n796 VSS.n783 147.374
R2466 VSS.n800 VSS.n784 147.374
R2467 VSS.n804 VSS.n785 147.374
R2468 VSS.n808 VSS.n786 147.374
R2469 VSS.n812 VSS.n787 147.374
R2470 VSS.n816 VSS.n788 147.374
R2471 VSS.n820 VSS.n789 147.374
R2472 VSS.n824 VSS.n790 147.374
R2473 VSS.n858 VSS.n791 147.374
R2474 VSS.n744 VSS.n683 147.374
R2475 VSS.n741 VSS.n684 147.374
R2476 VSS.n737 VSS.n685 147.374
R2477 VSS.n733 VSS.n686 147.374
R2478 VSS.n729 VSS.n687 147.374
R2479 VSS.n725 VSS.n688 147.374
R2480 VSS.n721 VSS.n689 147.374
R2481 VSS.n717 VSS.n690 147.374
R2482 VSS.n713 VSS.n691 147.374
R2483 VSS.n709 VSS.n692 147.374
R2484 VSS.n705 VSS.n693 147.374
R2485 VSS.n695 VSS.n693 147.374
R2486 VSS.n706 VSS.n692 147.374
R2487 VSS.n710 VSS.n691 147.374
R2488 VSS.n714 VSS.n690 147.374
R2489 VSS.n718 VSS.n689 147.374
R2490 VSS.n722 VSS.n688 147.374
R2491 VSS.n726 VSS.n687 147.374
R2492 VSS.n730 VSS.n686 147.374
R2493 VSS.n734 VSS.n685 147.374
R2494 VSS.n738 VSS.n684 147.374
R2495 VSS.n742 VSS.n683 147.374
R2496 VSS.n2123 VSS.n2122 147.374
R2497 VSS.n795 VSS.n782 147.374
R2498 VSS.n799 VSS.n783 147.374
R2499 VSS.n803 VSS.n784 147.374
R2500 VSS.n807 VSS.n785 147.374
R2501 VSS.n811 VSS.n786 147.374
R2502 VSS.n815 VSS.n787 147.374
R2503 VSS.n819 VSS.n788 147.374
R2504 VSS.n823 VSS.n789 147.374
R2505 VSS.n826 VSS.n790 147.374
R2506 VSS.n858 VSS.n857 147.374
R2507 VSS.n70 VSS.n46 140.69
R2508 VSS.n63 VSS.n46 140.69
R2509 VSS.n17 VSS.n16 140.69
R2510 VSS.n17 VSS.n8 140.69
R2511 VSS.n1276 VSS.n1275 140.69
R2512 VSS.n1275 VSS.n1249 140.69
R2513 VSS.n1268 VSS.n1249 140.69
R2514 VSS.n1268 VSS.n1267 140.69
R2515 VSS.n1267 VSS.n1253 140.69
R2516 VSS.n1260 VSS.n1253 140.69
R2517 VSS.n1260 VSS.n1259 140.69
R2518 VSS.n1209 VSS.n1204 140.69
R2519 VSS.n1216 VSS.n1204 140.69
R2520 VSS.n1217 VSS.n1216 140.69
R2521 VSS.n1217 VSS.n1200 140.69
R2522 VSS.n1225 VSS.n1200 140.69
R2523 VSS.n1226 VSS.n1225 140.69
R2524 VSS.n1226 VSS.n1197 140.69
R2525 VSS.n1354 VSS.n1348 140.69
R2526 VSS.n1355 VSS.n1354 140.69
R2527 VSS.n1355 VSS.n1344 140.69
R2528 VSS.n1362 VSS.n1344 140.69
R2529 VSS.n1363 VSS.n1362 140.69
R2530 VSS.n1363 VSS.n1340 140.69
R2531 VSS.n1370 VSS.n1340 140.69
R2532 VSS.n1871 VSS.n1839 140.69
R2533 VSS.n1864 VSS.n1839 140.69
R2534 VSS.n1864 VSS.n1863 140.69
R2535 VSS.n1863 VSS.n1843 140.69
R2536 VSS.n1856 VSS.n1843 140.69
R2537 VSS.n1856 VSS.n1855 140.69
R2538 VSS.n1855 VSS.n1847 140.69
R2539 VSS.n2254 VSS.n2253 117.233
R2540 VSS.n560 VSS.n543 99.5348
R2541 VSS.n566 VSS.n543 99.5348
R2542 VSS.n566 VSS.n539 99.5348
R2543 VSS.n573 VSS.n539 99.5348
R2544 VSS.n573 VSS.n535 99.5348
R2545 VSS.n579 VSS.n535 99.5348
R2546 VSS.n579 VSS.n443 99.5348
R2547 VSS.n2293 VSS.n445 99.5348
R2548 VSS.n2287 VSS.n445 99.5348
R2549 VSS.n2287 VSS.n2286 99.5348
R2550 VSS.n2286 VSS.n2285 99.5348
R2551 VSS.n2285 VSS.n454 99.5348
R2552 VSS.n2279 VSS.n454 99.5348
R2553 VSS.n2279 VSS.n2278 99.5348
R2554 VSS.n2278 VSS.n2277 99.5348
R2555 VSS.n2277 VSS.n461 99.5348
R2556 VSS.n2271 VSS.n461 99.5348
R2557 VSS.n2271 VSS.n2270 99.5348
R2558 VSS.n2270 VSS.n2269 99.5348
R2559 VSS.n2269 VSS.n468 99.5348
R2560 VSS.n2263 VSS.n468 99.5348
R2561 VSS.n2263 VSS.n2262 99.5348
R2562 VSS.n2262 VSS.n2261 99.5348
R2563 VSS.n2261 VSS.n475 99.5348
R2564 VSS.n2255 VSS.n475 99.5348
R2565 VSS.n2191 VSS.n654 99.5348
R2566 VSS.n2183 VSS.n2182 99.5348
R2567 VSS.n2182 VSS.n2181 99.5348
R2568 VSS.n2181 VSS.n662 99.5348
R2569 VSS.n1750 VSS.n671 99.5348
R2570 VSS.n2172 VSS.n671 99.5348
R2571 VSS.n2172 VSS.n2171 99.5348
R2572 VSS.n1307 VSS.n672 99.5348
R2573 VSS.n1308 VSS.n1307 99.5348
R2574 VSS.n1308 VSS.n681 99.5348
R2575 VSS.n1315 VSS.n682 99.5348
R2576 VSS.n1316 VSS.n1315 99.5348
R2577 VSS.n1323 VSS.n1322 99.5348
R2578 VSS.n1322 VSS.n1319 99.5348
R2579 VSS.n1922 VSS.n1921 99.5348
R2580 VSS.n1924 VSS.n1922 99.5348
R2581 VSS.n1924 VSS.n1923 99.5348
R2582 VSS.n1931 VSS.n1930 99.5348
R2583 VSS.n1932 VSS.n1931 99.5348
R2584 VSS.n1932 VSS.n859 99.5348
R2585 VSS.n1939 VSS.n860 99.5348
R2586 VSS.n1940 VSS.n1939 99.5348
R2587 VSS.n1940 VSS.n926 99.5348
R2588 VSS.n1956 VSS.n927 99.5348
R2589 VSS.n937 VSS.n927 99.5348
R2590 VSS.n938 VSS.n937 99.5348
R2591 VSS.n1175 VSS.n1174 99.5348
R2592 VSS.t0 VSS.n654 92.2161
R2593 VSS.n1175 VSS.t40 92.2161
R2594 VSS.n321 VSS.t81 90.6265
R2595 VSS.n305 VSS.t74 90.6265
R2596 VSS.n377 VSS.t90 90.6265
R2597 VSS.n360 VSS.t84 90.6265
R2598 VSS.t5 VSS.n1323 89.2886
R2599 VSS.n1319 VSS.t23 89.2886
R2600 VSS.n562 VSS.n545 85.8358
R2601 VSS.n558 VSS.n557 85.8358
R2602 VSS.n641 VSS.n640 85.8358
R2603 VSS.n1721 VSS.n1720 82.4476
R2604 VSS.n1810 VSS.n1809 82.4476
R2605 VSS.n1682 VSS.n1679 82.4476
R2606 VSS.n2011 VSS.n876 82.4476
R2607 VSS.n2083 VSS.n2082 82.4476
R2608 VSS.n2017 VSS.n924 82.4476
R2609 VSS.n2038 VSS.n2035 82.4476
R2610 VSS.n746 VSS.n745 82.4476
R2611 VSS.n2160 VSS.n2159 82.4476
R2612 VSS.n2126 VSS.n2125 82.4476
R2613 VSS.n856 VSS.n855 82.4476
R2614 VSS.n321 VSS.t79 81.8918
R2615 VSS.n320 VSS.t121 81.8918
R2616 VSS.n305 VSS.t71 81.8918
R2617 VSS.n381 VSS.t87 81.8918
R2618 VSS.n377 VSS.t89 81.8918
R2619 VSS.n360 VSS.t82 81.8918
R2620 VSS.n48 VSS.t85 81.8918
R2621 VSS.n61 VSS.t108 81.8918
R2622 VSS.n7 VSS.t119 81.8918
R2623 VSS.n24 VSS.t117 81.8918
R2624 VSS.n1316 VSS.n701 79.0424
R2625 VSS.n433 VSS.n218 76.8005
R2626 VSS.n2553 VSS.n2498 76.8005
R2627 VSS.n429 VSS.n428 76.8005
R2628 VSS.n2492 VSS.n2491 76.8005
R2629 VSS.n1170 VSS.n952 76.8005
R2630 VSS.n2097 VSS.n886 76.8005
R2631 VSS.n1728 VSS.n1727 76.8005
R2632 VSS.n2189 VSS.n657 76.8005
R2633 VSS.n2295 VSS.n443 74.6512
R2634 VSS.t22 VSS.n662 71.7237
R2635 VSS.t18 VSS.n1956 71.7237
R2636 VSS.n63 VSS.t110 70.3453
R2637 VSS.t120 VSS.n8 70.3453
R2638 VSS.n1259 VSS.t105 70.3453
R2639 VSS.t63 VSS.n1197 70.3453
R2640 VSS.t68 VSS.n1348 70.3453
R2641 VSS.t70 VSS.n1871 70.3453
R2642 VSS.t15 VSS.n682 68.7962
R2643 VSS.n1923 VSS.t41 68.7962
R2644 VSS.n2079 VSS.n899 66.162
R2645 VSS.n1129 VSS.n1128 64.7534
R2646 VSS.n1517 VSS.n1516 64.7534
R2647 VSS.n2202 VSS.n2201 62.1181
R2648 VSS.n1724 VSS.n98 61.9943
R2649 VSS.n431 VSS.n220 54.18
R2650 VSS.n2556 VSS.n80 54.18
R2651 VSS.n2171 VSS.t16 51.2314
R2652 VSS.t17 VSS.n860 51.2314
R2653 VSS.n2255 VSS.t32 49.7676
R2654 VSS.t16 VSS.n672 48.3039
R2655 VSS.t17 VSS.n859 48.3039
R2656 VSS.n1764 VSS.n1763 45.3391
R2657 VSS.n1081 VSS.n1080 39.1534
R2658 VSS.n1033 VSS.n1032 39.1534
R2659 VSS.n1565 VSS.n1564 39.1534
R2660 VSS.n1613 VSS.n1612 39.1534
R2661 VSS.t32 VSS.n2254 38.2032
R2662 VSS.n431 VSS.n216 35.4256
R2663 VSS.n437 VSS.n216 35.4256
R2664 VSS.n2296 VSS.n212 35.4256
R2665 VSS.n2302 VSS.n205 35.4256
R2666 VSS.n2309 VSS.n205 35.4256
R2667 VSS.n2309 VSS.n2308 35.4256
R2668 VSS.n2315 VSS.n198 35.4256
R2669 VSS.n2322 VSS.n198 35.4256
R2670 VSS.n2322 VSS.n2321 35.4256
R2671 VSS.n2328 VSS.n191 35.4256
R2672 VSS.n2335 VSS.n191 35.4256
R2673 VSS.n2335 VSS.n2334 35.4256
R2674 VSS.n2341 VSS.n184 35.4256
R2675 VSS.n2348 VSS.n184 35.4256
R2676 VSS.n2348 VSS.n2347 35.4256
R2677 VSS.n2354 VSS.n177 35.4256
R2678 VSS.n2360 VSS.n177 35.4256
R2679 VSS.n2366 VSS.n173 35.4256
R2680 VSS.n2366 VSS.n169 35.4256
R2681 VSS.n2372 VSS.n169 35.4256
R2682 VSS.n2378 VSS.n165 35.4256
R2683 VSS.n2378 VSS.n161 35.4256
R2684 VSS.n2384 VSS.n161 35.4256
R2685 VSS.n2390 VSS.n157 35.4256
R2686 VSS.n2390 VSS.n153 35.4256
R2687 VSS.n2396 VSS.n153 35.4256
R2688 VSS.n2402 VSS.n148 35.4256
R2689 VSS.n2402 VSS.n149 35.4256
R2690 VSS.n2408 VSS.n140 35.4256
R2691 VSS.n2414 VSS.n140 35.4256
R2692 VSS.n2414 VSS.n141 35.4256
R2693 VSS.n2420 VSS.n132 35.4256
R2694 VSS.n2426 VSS.n132 35.4256
R2695 VSS.n2426 VSS.n133 35.4256
R2696 VSS.n2432 VSS.n124 35.4256
R2697 VSS.n2438 VSS.n124 35.4256
R2698 VSS.n2438 VSS.n125 35.4256
R2699 VSS.n2444 VSS.n116 35.4256
R2700 VSS.n2450 VSS.n116 35.4256
R2701 VSS.n2450 VSS.n117 35.4256
R2702 VSS.n2456 VSS.n109 35.4256
R2703 VSS.n2462 VSS.n109 35.4256
R2704 VSS.n2495 VSS.n104 35.4256
R2705 VSS.n2495 VSS.n80 35.4256
R2706 VSS.n1723 VSS.n1657 35.4256
R2707 VSS.n2170 VSS.n674 35.4256
R2708 VSS.n2164 VSS.n2163 35.4256
R2709 VSS.n1329 VSS.n694 35.4256
R2710 VSS.n781 VSS.n775 35.4256
R2711 VSS.n2120 VSS.n861 35.4256
R2712 VSS.n1959 VSS.n1957 35.4256
R2713 VSS.n2094 VSS.n890 35.4256
R2714 VSS.n2088 VSS.n890 35.4256
R2715 VSS.n2088 VSS.n2087 35.4256
R2716 VSS.n2086 VSS.n899 35.4256
R2717 VSS.n2354 VSS.t7 34.9046
R2718 VSS.n149 VSS.t11 34.9046
R2719 VSS.t83 VSS.n212 33.8627
R2720 VSS.n2462 VSS.t72 33.8627
R2721 VSS.n312 VSS.n311 32.8962
R2722 VSS.n367 VSS.n366 32.8962
R2723 VSS.t15 VSS.n681 30.739
R2724 VSS.n1930 VSS.t41 30.739
R2725 VSS.n2295 VSS.n2294 30.7369
R2726 VSS.n2294 VSS.t52 29.695
R2727 VSS.n2456 VSS.t36 29.695
R2728 VSS.n2360 VSS.t13 28.6531
R2729 VSS.t45 VSS.n148 28.6531
R2730 VSS.n64 VSS.n62 28.3989
R2731 VSS.n21 VSS.n20 28.3989
R2732 VSS.n336 VSS.n335 27.9576
R2733 VSS.n340 VSS.n339 27.9576
R2734 VSS.n344 VSS.n343 27.9576
R2735 VSS.n348 VSS.n347 27.9576
R2736 VSS.n352 VSS.n351 27.9576
R2737 VSS.t22 VSS.n1750 27.8115
R2738 VSS.t18 VSS.n926 27.8115
R2739 VSS.n334 VSS.n333 27.7293
R2740 VSS.n338 VSS.n337 27.7293
R2741 VSS.n342 VSS.n341 27.7293
R2742 VSS.n346 VSS.n345 27.7293
R2743 VSS.n350 VSS.n349 27.7293
R2744 VSS.n354 VSS.n353 27.7293
R2745 VSS.n42 VSS.n41 27.7293
R2746 VSS.n40 VSS.n39 27.7293
R2747 VSS.n38 VSS.n37 27.7293
R2748 VSS.n36 VSS.n35 27.7293
R2749 VSS.n34 VSS.n33 27.7293
R2750 VSS.n2341 VSS.t30 27.6112
R2751 VSS.n141 VSS.t1 27.6112
R2752 VSS.n2013 VSS.n861 27.6112
R2753 VSS.n328 VSS.n299 27.5286
R2754 VSS.n329 VSS.n297 27.5286
R2755 VSS.n389 VSS.n372 27.5286
R2756 VSS.n388 VSS.n374 27.5286
R2757 VSS.n58 VSS.n49 27.5286
R2758 VSS.n29 VSS.n6 27.5286
R2759 VSS.n1280 VSS.n1246 25.6009
R2760 VSS.n1208 VSS.n1196 25.6009
R2761 VSS.n1372 VSS.n1371 25.6009
R2762 VSS.n1849 VSS.n1386 25.6009
R2763 VSS.n434 VSS.n433 25.6005
R2764 VSS.n435 VSS.n434 25.6005
R2765 VSS.n435 VSS.n210 25.6005
R2766 VSS.n2298 VSS.n210 25.6005
R2767 VSS.n2299 VSS.n2298 25.6005
R2768 VSS.n2300 VSS.n2299 25.6005
R2769 VSS.n2300 VSS.n203 25.6005
R2770 VSS.n2311 VSS.n203 25.6005
R2771 VSS.n2312 VSS.n2311 25.6005
R2772 VSS.n2313 VSS.n2312 25.6005
R2773 VSS.n2313 VSS.n196 25.6005
R2774 VSS.n2324 VSS.n196 25.6005
R2775 VSS.n2325 VSS.n2324 25.6005
R2776 VSS.n2326 VSS.n2325 25.6005
R2777 VSS.n2326 VSS.n189 25.6005
R2778 VSS.n2337 VSS.n189 25.6005
R2779 VSS.n2338 VSS.n2337 25.6005
R2780 VSS.n2339 VSS.n2338 25.6005
R2781 VSS.n2339 VSS.n182 25.6005
R2782 VSS.n2350 VSS.n182 25.6005
R2783 VSS.n2351 VSS.n2350 25.6005
R2784 VSS.n2352 VSS.n2351 25.6005
R2785 VSS.n2352 VSS.n175 25.6005
R2786 VSS.n2362 VSS.n175 25.6005
R2787 VSS.n2363 VSS.n2362 25.6005
R2788 VSS.n2364 VSS.n2363 25.6005
R2789 VSS.n2364 VSS.n167 25.6005
R2790 VSS.n2374 VSS.n167 25.6005
R2791 VSS.n2375 VSS.n2374 25.6005
R2792 VSS.n2376 VSS.n2375 25.6005
R2793 VSS.n2376 VSS.n159 25.6005
R2794 VSS.n2386 VSS.n159 25.6005
R2795 VSS.n2387 VSS.n2386 25.6005
R2796 VSS.n2388 VSS.n2387 25.6005
R2797 VSS.n2388 VSS.n151 25.6005
R2798 VSS.n2398 VSS.n151 25.6005
R2799 VSS.n2399 VSS.n2398 25.6005
R2800 VSS.n2400 VSS.n2399 25.6005
R2801 VSS.n2400 VSS.n143 25.6005
R2802 VSS.n2410 VSS.n143 25.6005
R2803 VSS.n2411 VSS.n2410 25.6005
R2804 VSS.n2412 VSS.n2411 25.6005
R2805 VSS.n2412 VSS.n135 25.6005
R2806 VSS.n2422 VSS.n135 25.6005
R2807 VSS.n2423 VSS.n2422 25.6005
R2808 VSS.n2424 VSS.n2423 25.6005
R2809 VSS.n2424 VSS.n127 25.6005
R2810 VSS.n2434 VSS.n127 25.6005
R2811 VSS.n2435 VSS.n2434 25.6005
R2812 VSS.n2436 VSS.n2435 25.6005
R2813 VSS.n2436 VSS.n119 25.6005
R2814 VSS.n2446 VSS.n119 25.6005
R2815 VSS.n2447 VSS.n2446 25.6005
R2816 VSS.n2448 VSS.n2447 25.6005
R2817 VSS.n2448 VSS.n111 25.6005
R2818 VSS.n2458 VSS.n111 25.6005
R2819 VSS.n2459 VSS.n2458 25.6005
R2820 VSS.n2460 VSS.n2459 25.6005
R2821 VSS.n2460 VSS.n102 25.6005
R2822 VSS.n2497 VSS.n102 25.6005
R2823 VSS.n2498 VSS.n2497 25.6005
R2824 VSS.n246 VSS.n218 25.6005
R2825 VSS.n247 VSS.n246 25.6005
R2826 VSS.n248 VSS.n247 25.6005
R2827 VSS.n248 VSS.n242 25.6005
R2828 VSS.n254 VSS.n242 25.6005
R2829 VSS.n255 VSS.n254 25.6005
R2830 VSS.n256 VSS.n255 25.6005
R2831 VSS.n256 VSS.n240 25.6005
R2832 VSS.n262 VSS.n240 25.6005
R2833 VSS.n263 VSS.n262 25.6005
R2834 VSS.n264 VSS.n263 25.6005
R2835 VSS.n264 VSS.n238 25.6005
R2836 VSS.n270 VSS.n238 25.6005
R2837 VSS.n271 VSS.n270 25.6005
R2838 VSS.n280 VSS.n234 25.6005
R2839 VSS.n292 VSS.n232 25.6005
R2840 VSS.n397 VSS.n228 25.6005
R2841 VSS.n403 VSS.n228 25.6005
R2842 VSS.n404 VSS.n403 25.6005
R2843 VSS.n405 VSS.n404 25.6005
R2844 VSS.n405 VSS.n226 25.6005
R2845 VSS.n411 VSS.n226 25.6005
R2846 VSS.n412 VSS.n411 25.6005
R2847 VSS.n413 VSS.n412 25.6005
R2848 VSS.n413 VSS.n224 25.6005
R2849 VSS.n419 VSS.n224 25.6005
R2850 VSS.n420 VSS.n419 25.6005
R2851 VSS.n421 VSS.n420 25.6005
R2852 VSS.n421 VSS.n222 25.6005
R2853 VSS.n427 VSS.n222 25.6005
R2854 VSS.n428 VSS.n427 25.6005
R2855 VSS.n429 VSS.n214 25.6005
R2856 VSS.n439 VSS.n214 25.6005
R2857 VSS.n440 VSS.n439 25.6005
R2858 VSS.n441 VSS.n440 25.6005
R2859 VSS.n441 VSS.n207 25.6005
R2860 VSS.n2304 VSS.n207 25.6005
R2861 VSS.n2305 VSS.n2304 25.6005
R2862 VSS.n2306 VSS.n2305 25.6005
R2863 VSS.n2306 VSS.n200 25.6005
R2864 VSS.n2317 VSS.n200 25.6005
R2865 VSS.n2318 VSS.n2317 25.6005
R2866 VSS.n2319 VSS.n2318 25.6005
R2867 VSS.n2319 VSS.n193 25.6005
R2868 VSS.n2330 VSS.n193 25.6005
R2869 VSS.n2331 VSS.n2330 25.6005
R2870 VSS.n2332 VSS.n2331 25.6005
R2871 VSS.n2332 VSS.n186 25.6005
R2872 VSS.n2343 VSS.n186 25.6005
R2873 VSS.n2344 VSS.n2343 25.6005
R2874 VSS.n2345 VSS.n2344 25.6005
R2875 VSS.n2345 VSS.n179 25.6005
R2876 VSS.n2356 VSS.n179 25.6005
R2877 VSS.n2357 VSS.n2356 25.6005
R2878 VSS.n2358 VSS.n2357 25.6005
R2879 VSS.n2358 VSS.n171 25.6005
R2880 VSS.n2368 VSS.n171 25.6005
R2881 VSS.n2369 VSS.n2368 25.6005
R2882 VSS.n2370 VSS.n2369 25.6005
R2883 VSS.n2370 VSS.n163 25.6005
R2884 VSS.n2380 VSS.n163 25.6005
R2885 VSS.n2381 VSS.n2380 25.6005
R2886 VSS.n2382 VSS.n2381 25.6005
R2887 VSS.n2382 VSS.n155 25.6005
R2888 VSS.n2392 VSS.n155 25.6005
R2889 VSS.n2393 VSS.n2392 25.6005
R2890 VSS.n2394 VSS.n2393 25.6005
R2891 VSS.n2394 VSS.n146 25.6005
R2892 VSS.n2404 VSS.n146 25.6005
R2893 VSS.n2405 VSS.n2404 25.6005
R2894 VSS.n2406 VSS.n2405 25.6005
R2895 VSS.n2406 VSS.n138 25.6005
R2896 VSS.n2416 VSS.n138 25.6005
R2897 VSS.n2417 VSS.n2416 25.6005
R2898 VSS.n2418 VSS.n2417 25.6005
R2899 VSS.n2418 VSS.n130 25.6005
R2900 VSS.n2428 VSS.n130 25.6005
R2901 VSS.n2429 VSS.n2428 25.6005
R2902 VSS.n2430 VSS.n2429 25.6005
R2903 VSS.n2430 VSS.n122 25.6005
R2904 VSS.n2440 VSS.n122 25.6005
R2905 VSS.n2441 VSS.n2440 25.6005
R2906 VSS.n2442 VSS.n2441 25.6005
R2907 VSS.n2442 VSS.n114 25.6005
R2908 VSS.n2452 VSS.n114 25.6005
R2909 VSS.n2453 VSS.n2452 25.6005
R2910 VSS.n2454 VSS.n2453 25.6005
R2911 VSS.n2454 VSS.n107 25.6005
R2912 VSS.n2464 VSS.n107 25.6005
R2913 VSS.n2465 VSS.n2464 25.6005
R2914 VSS.n2493 VSS.n2465 25.6005
R2915 VSS.n2493 VSS.n2492 25.6005
R2916 VSS.n2553 VSS.n2552 25.6005
R2917 VSS.n2552 VSS.n2551 25.6005
R2918 VSS.n2551 VSS.n2550 25.6005
R2919 VSS.n2550 VSS.n2548 25.6005
R2920 VSS.n2548 VSS.n2545 25.6005
R2921 VSS.n2545 VSS.n2544 25.6005
R2922 VSS.n2544 VSS.n2541 25.6005
R2923 VSS.n2541 VSS.n2540 25.6005
R2924 VSS.n2540 VSS.n2537 25.6005
R2925 VSS.n2537 VSS.n2536 25.6005
R2926 VSS.n2536 VSS.n2533 25.6005
R2927 VSS.n2533 VSS.n2532 25.6005
R2928 VSS.n2532 VSS.n2529 25.6005
R2929 VSS.n2529 VSS.n2528 25.6005
R2930 VSS.n2520 VSS.n2517 25.6005
R2931 VSS.n2506 VSS.n2503 25.6005
R2932 VSS.n2559 VSS.n76 25.6005
R2933 VSS.n2559 VSS.n77 25.6005
R2934 VSS.n2466 VSS.n77 25.6005
R2935 VSS.n2469 VSS.n2466 25.6005
R2936 VSS.n2470 VSS.n2469 25.6005
R2937 VSS.n2473 VSS.n2470 25.6005
R2938 VSS.n2474 VSS.n2473 25.6005
R2939 VSS.n2477 VSS.n2474 25.6005
R2940 VSS.n2478 VSS.n2477 25.6005
R2941 VSS.n2481 VSS.n2478 25.6005
R2942 VSS.n2482 VSS.n2481 25.6005
R2943 VSS.n2485 VSS.n2482 25.6005
R2944 VSS.n2486 VSS.n2485 25.6005
R2945 VSS.n2489 VSS.n2486 25.6005
R2946 VSS.n2491 VSS.n2489 25.6005
R2947 VSS.n1721 VSS.n1429 25.6005
R2948 VSS.n1738 VSS.n1429 25.6005
R2949 VSS.n1739 VSS.n1738 25.6005
R2950 VSS.n1740 VSS.n1739 25.6005
R2951 VSS.n1740 VSS.n1401 25.6005
R2952 VSS.n1829 VSS.n1401 25.6005
R2953 VSS.n1829 VSS.n1828 25.6005
R2954 VSS.n1828 VSS.n1827 25.6005
R2955 VSS.n1827 VSS.n1402 25.6005
R2956 VSS.n1811 VSS.n1402 25.6005
R2957 VSS.n1811 VSS.n1810 25.6005
R2958 VSS.n1720 VSS.n1719 25.6005
R2959 VSS.n1719 VSS.n1659 25.6005
R2960 VSS.n1660 VSS.n1659 25.6005
R2961 VSS.n1712 VSS.n1660 25.6005
R2962 VSS.n1712 VSS.n1711 25.6005
R2963 VSS.n1711 VSS.n1710 25.6005
R2964 VSS.n1710 VSS.n1662 25.6005
R2965 VSS.n1705 VSS.n1662 25.6005
R2966 VSS.n1705 VSS.n1704 25.6005
R2967 VSS.n1704 VSS.n1703 25.6005
R2968 VSS.n1703 VSS.n1665 25.6005
R2969 VSS.n1698 VSS.n1665 25.6005
R2970 VSS.n1698 VSS.n1697 25.6005
R2971 VSS.n1697 VSS.n1696 25.6005
R2972 VSS.n1696 VSS.n1668 25.6005
R2973 VSS.n1691 VSS.n1668 25.6005
R2974 VSS.n1691 VSS.n1690 25.6005
R2975 VSS.n1690 VSS.n1689 25.6005
R2976 VSS.n1689 VSS.n1671 25.6005
R2977 VSS.n1684 VSS.n1671 25.6005
R2978 VSS.n1684 VSS.n1683 25.6005
R2979 VSS.n1683 VSS.n1682 25.6005
R2980 VSS.n1679 VSS.n1678 25.6005
R2981 VSS.n1678 VSS.n1676 25.6005
R2982 VSS.n1676 VSS.n1675 25.6005
R2983 VSS.n1675 VSS.n1425 25.6005
R2984 VSS.n1746 VSS.n1425 25.6005
R2985 VSS.n1747 VSS.n1746 25.6005
R2986 VSS.n1760 VSS.n1759 25.6005
R2987 VSS.n1809 VSS.n1411 25.6005
R2988 VSS.n1804 VSS.n1411 25.6005
R2989 VSS.n1804 VSS.n1803 25.6005
R2990 VSS.n1803 VSS.n1802 25.6005
R2991 VSS.n1802 VSS.n1413 25.6005
R2992 VSS.n1796 VSS.n1413 25.6005
R2993 VSS.n1796 VSS.n1795 25.6005
R2994 VSS.n1795 VSS.n1794 25.6005
R2995 VSS.n1794 VSS.n1415 25.6005
R2996 VSS.n1788 VSS.n1415 25.6005
R2997 VSS.n1788 VSS.n1787 25.6005
R2998 VSS.n1787 VSS.n1786 25.6005
R2999 VSS.n1786 VSS.n1417 25.6005
R3000 VSS.n1780 VSS.n1417 25.6005
R3001 VSS.n1780 VSS.n1779 25.6005
R3002 VSS.n1779 VSS.n1778 25.6005
R3003 VSS.n1778 VSS.n1419 25.6005
R3004 VSS.n1772 VSS.n1419 25.6005
R3005 VSS.n1772 VSS.n1771 25.6005
R3006 VSS.n1771 VSS.n1770 25.6005
R3007 VSS.n1770 VSS.n1421 25.6005
R3008 VSS.n1764 VSS.n1421 25.6005
R3009 VSS.n1170 VSS.n1169 25.6005
R3010 VSS.n1169 VSS.n1168 25.6005
R3011 VSS.n1168 VSS.n1167 25.6005
R3012 VSS.n1167 VSS.n1165 25.6005
R3013 VSS.n1165 VSS.n1162 25.6005
R3014 VSS.n1162 VSS.n1161 25.6005
R3015 VSS.n1161 VSS.n1158 25.6005
R3016 VSS.n1158 VSS.n1157 25.6005
R3017 VSS.n1157 VSS.n1154 25.6005
R3018 VSS.n1154 VSS.n1153 25.6005
R3019 VSS.n1153 VSS.n1150 25.6005
R3020 VSS.n1150 VSS.n1149 25.6005
R3021 VSS.n1149 VSS.n1146 25.6005
R3022 VSS.n1146 VSS.n1145 25.6005
R3023 VSS.n1145 VSS.n1142 25.6005
R3024 VSS.n1142 VSS.n1141 25.6005
R3025 VSS.n1141 VSS.n1138 25.6005
R3026 VSS.n1138 VSS.n1137 25.6005
R3027 VSS.n1137 VSS.n1135 25.6005
R3028 VSS.n1135 VSS.n1134 25.6005
R3029 VSS.n1134 VSS.n953 25.6005
R3030 VSS.n1129 VSS.n953 25.6005
R3031 VSS.n1128 VSS.n1127 25.6005
R3032 VSS.n1127 VSS.n955 25.6005
R3033 VSS.n1121 VSS.n955 25.6005
R3034 VSS.n1121 VSS.n1120 25.6005
R3035 VSS.n1120 VSS.n1119 25.6005
R3036 VSS.n1119 VSS.n957 25.6005
R3037 VSS.n1113 VSS.n957 25.6005
R3038 VSS.n1113 VSS.n1112 25.6005
R3039 VSS.n1112 VSS.n1111 25.6005
R3040 VSS.n1111 VSS.n959 25.6005
R3041 VSS.n1105 VSS.n959 25.6005
R3042 VSS.n1105 VSS.n1104 25.6005
R3043 VSS.n1104 VSS.n1103 25.6005
R3044 VSS.n1103 VSS.n961 25.6005
R3045 VSS.n1097 VSS.n961 25.6005
R3046 VSS.n1097 VSS.n1096 25.6005
R3047 VSS.n1096 VSS.n1095 25.6005
R3048 VSS.n1095 VSS.n963 25.6005
R3049 VSS.n1089 VSS.n963 25.6005
R3050 VSS.n1089 VSS.n1088 25.6005
R3051 VSS.n1088 VSS.n1087 25.6005
R3052 VSS.n1087 VSS.n965 25.6005
R3053 VSS.n1081 VSS.n965 25.6005
R3054 VSS.n1080 VSS.n1079 25.6005
R3055 VSS.n1079 VSS.n967 25.6005
R3056 VSS.n1073 VSS.n967 25.6005
R3057 VSS.n1073 VSS.n1072 25.6005
R3058 VSS.n1072 VSS.n1071 25.6005
R3059 VSS.n1071 VSS.n969 25.6005
R3060 VSS.n1065 VSS.n969 25.6005
R3061 VSS.n1065 VSS.n1064 25.6005
R3062 VSS.n1064 VSS.n1063 25.6005
R3063 VSS.n1063 VSS.n971 25.6005
R3064 VSS.n1057 VSS.n971 25.6005
R3065 VSS.n1057 VSS.n1056 25.6005
R3066 VSS.n1056 VSS.n1055 25.6005
R3067 VSS.n1055 VSS.n973 25.6005
R3068 VSS.n1049 VSS.n973 25.6005
R3069 VSS.n1049 VSS.n1048 25.6005
R3070 VSS.n1048 VSS.n1047 25.6005
R3071 VSS.n1047 VSS.n975 25.6005
R3072 VSS.n1041 VSS.n975 25.6005
R3073 VSS.n1041 VSS.n1040 25.6005
R3074 VSS.n1040 VSS.n1039 25.6005
R3075 VSS.n1039 VSS.n977 25.6005
R3076 VSS.n1033 VSS.n977 25.6005
R3077 VSS.n1032 VSS.n1031 25.6005
R3078 VSS.n1031 VSS.n979 25.6005
R3079 VSS.n1025 VSS.n979 25.6005
R3080 VSS.n1025 VSS.n1024 25.6005
R3081 VSS.n1024 VSS.n1023 25.6005
R3082 VSS.n1023 VSS.n981 25.6005
R3083 VSS.n1017 VSS.n981 25.6005
R3084 VSS.n1017 VSS.n1016 25.6005
R3085 VSS.n1016 VSS.n1015 25.6005
R3086 VSS.n1015 VSS.n983 25.6005
R3087 VSS.n1009 VSS.n983 25.6005
R3088 VSS.n1009 VSS.n1008 25.6005
R3089 VSS.n1008 VSS.n1007 25.6005
R3090 VSS.n1007 VSS.n985 25.6005
R3091 VSS.n1001 VSS.n985 25.6005
R3092 VSS.n1001 VSS.n1000 25.6005
R3093 VSS.n1000 VSS.n999 25.6005
R3094 VSS.n999 VSS.n987 25.6005
R3095 VSS.n993 VSS.n987 25.6005
R3096 VSS.n993 VSS.n992 25.6005
R3097 VSS.n992 VSS.n991 25.6005
R3098 VSS.n991 VSS.n886 25.6005
R3099 VSS.n1730 VSS.n1393 25.6005
R3100 VSS.n1834 VSS.n1394 25.6005
R3101 VSS.n1822 VSS.n1816 25.6005
R3102 VSS.n1817 VSS.n677 25.6005
R3103 VSS.n2168 VSS.n677 25.6005
R3104 VSS.n2168 VSS.n2167 25.6005
R3105 VSS.n2167 VSS.n2166 25.6005
R3106 VSS.n2166 VSS.n678 25.6005
R3107 VSS.n1326 VSS.n678 25.6005
R3108 VSS.n1331 VSS.n1326 25.6005
R3109 VSS.n1902 VSS.n754 25.6005
R3110 VSS.n2147 VSS.n754 25.6005
R3111 VSS.n2147 VSS.n2146 25.6005
R3112 VSS.n2146 VSS.n2145 25.6005
R3113 VSS.n2133 VSS.n770 25.6005
R3114 VSS.n2133 VSS.n2132 25.6005
R3115 VSS.n2132 VSS.n2131 25.6005
R3116 VSS.n2131 VSS.n771 25.6005
R3117 VSS.n864 VSS.n771 25.6005
R3118 VSS.n2118 VSS.n864 25.6005
R3119 VSS.n2118 VSS.n2117 25.6005
R3120 VSS.n867 VSS.n865 25.6005
R3121 VSS.n2113 VSS.n868 25.6005
R3122 VSS.n2101 VSS.n883 25.6005
R3123 VSS.n1473 VSS.n657 25.6005
R3124 VSS.n1476 VSS.n1473 25.6005
R3125 VSS.n1477 VSS.n1476 25.6005
R3126 VSS.n1480 VSS.n1477 25.6005
R3127 VSS.n1481 VSS.n1480 25.6005
R3128 VSS.n1484 VSS.n1481 25.6005
R3129 VSS.n1485 VSS.n1484 25.6005
R3130 VSS.n1488 VSS.n1485 25.6005
R3131 VSS.n1489 VSS.n1488 25.6005
R3132 VSS.n1492 VSS.n1489 25.6005
R3133 VSS.n1493 VSS.n1492 25.6005
R3134 VSS.n1496 VSS.n1493 25.6005
R3135 VSS.n1497 VSS.n1496 25.6005
R3136 VSS.n1500 VSS.n1497 25.6005
R3137 VSS.n1501 VSS.n1500 25.6005
R3138 VSS.n1504 VSS.n1501 25.6005
R3139 VSS.n1505 VSS.n1504 25.6005
R3140 VSS.n1508 VSS.n1505 25.6005
R3141 VSS.n1509 VSS.n1508 25.6005
R3142 VSS.n1512 VSS.n1509 25.6005
R3143 VSS.n1513 VSS.n1512 25.6005
R3144 VSS.n1516 VSS.n1513 25.6005
R3145 VSS.n1520 VSS.n1517 25.6005
R3146 VSS.n1521 VSS.n1520 25.6005
R3147 VSS.n1524 VSS.n1521 25.6005
R3148 VSS.n1525 VSS.n1524 25.6005
R3149 VSS.n1528 VSS.n1525 25.6005
R3150 VSS.n1529 VSS.n1528 25.6005
R3151 VSS.n1532 VSS.n1529 25.6005
R3152 VSS.n1533 VSS.n1532 25.6005
R3153 VSS.n1536 VSS.n1533 25.6005
R3154 VSS.n1537 VSS.n1536 25.6005
R3155 VSS.n1540 VSS.n1537 25.6005
R3156 VSS.n1541 VSS.n1540 25.6005
R3157 VSS.n1544 VSS.n1541 25.6005
R3158 VSS.n1545 VSS.n1544 25.6005
R3159 VSS.n1548 VSS.n1545 25.6005
R3160 VSS.n1549 VSS.n1548 25.6005
R3161 VSS.n1552 VSS.n1549 25.6005
R3162 VSS.n1553 VSS.n1552 25.6005
R3163 VSS.n1556 VSS.n1553 25.6005
R3164 VSS.n1557 VSS.n1556 25.6005
R3165 VSS.n1560 VSS.n1557 25.6005
R3166 VSS.n1561 VSS.n1560 25.6005
R3167 VSS.n1564 VSS.n1561 25.6005
R3168 VSS.n1568 VSS.n1565 25.6005
R3169 VSS.n1569 VSS.n1568 25.6005
R3170 VSS.n1572 VSS.n1569 25.6005
R3171 VSS.n1573 VSS.n1572 25.6005
R3172 VSS.n1576 VSS.n1573 25.6005
R3173 VSS.n1577 VSS.n1576 25.6005
R3174 VSS.n1580 VSS.n1577 25.6005
R3175 VSS.n1581 VSS.n1580 25.6005
R3176 VSS.n1584 VSS.n1581 25.6005
R3177 VSS.n1585 VSS.n1584 25.6005
R3178 VSS.n1588 VSS.n1585 25.6005
R3179 VSS.n1589 VSS.n1588 25.6005
R3180 VSS.n1592 VSS.n1589 25.6005
R3181 VSS.n1593 VSS.n1592 25.6005
R3182 VSS.n1596 VSS.n1593 25.6005
R3183 VSS.n1597 VSS.n1596 25.6005
R3184 VSS.n1600 VSS.n1597 25.6005
R3185 VSS.n1601 VSS.n1600 25.6005
R3186 VSS.n1604 VSS.n1601 25.6005
R3187 VSS.n1605 VSS.n1604 25.6005
R3188 VSS.n1608 VSS.n1605 25.6005
R3189 VSS.n1609 VSS.n1608 25.6005
R3190 VSS.n1612 VSS.n1609 25.6005
R3191 VSS.n1616 VSS.n1613 25.6005
R3192 VSS.n1617 VSS.n1616 25.6005
R3193 VSS.n1620 VSS.n1617 25.6005
R3194 VSS.n1621 VSS.n1620 25.6005
R3195 VSS.n1624 VSS.n1621 25.6005
R3196 VSS.n1625 VSS.n1624 25.6005
R3197 VSS.n1628 VSS.n1625 25.6005
R3198 VSS.n1629 VSS.n1628 25.6005
R3199 VSS.n1632 VSS.n1629 25.6005
R3200 VSS.n1633 VSS.n1632 25.6005
R3201 VSS.n1636 VSS.n1633 25.6005
R3202 VSS.n1637 VSS.n1636 25.6005
R3203 VSS.n1640 VSS.n1637 25.6005
R3204 VSS.n1641 VSS.n1640 25.6005
R3205 VSS.n1644 VSS.n1641 25.6005
R3206 VSS.n1645 VSS.n1644 25.6005
R3207 VSS.n1648 VSS.n1645 25.6005
R3208 VSS.n1650 VSS.n1648 25.6005
R3209 VSS.n1651 VSS.n1650 25.6005
R3210 VSS.n1652 VSS.n1651 25.6005
R3211 VSS.n1652 VSS.n1435 25.6005
R3212 VSS.n1727 VSS.n1435 25.6005
R3213 VSS.n2185 VSS.n660 25.6005
R3214 VSS.n2179 VSS.n2178 25.6005
R3215 VSS.n667 VSS.n665 25.6005
R3216 VSS.n2174 VSS.n668 25.6005
R3217 VSS.n1304 VSS.n668 25.6005
R3218 VSS.n1305 VSS.n1304 25.6005
R3219 VSS.n1305 VSS.n1302 25.6005
R3220 VSS.n1311 VSS.n1302 25.6005
R3221 VSS.n1312 VSS.n1311 25.6005
R3222 VSS.n1313 VSS.n1312 25.6005
R3223 VSS.n1908 VSS.n1300 25.6005
R3224 VSS.n1320 VSS.n1300 25.6005
R3225 VSS.n1320 VSS.n1192 25.6005
R3226 VSS.n1919 VSS.n1192 25.6005
R3227 VSS.n1927 VSS.n1926 25.6005
R3228 VSS.n1928 VSS.n1927 25.6005
R3229 VSS.n1928 VSS.n1185 25.6005
R3230 VSS.n1934 VSS.n1185 25.6005
R3231 VSS.n1935 VSS.n1934 25.6005
R3232 VSS.n1936 VSS.n1935 25.6005
R3233 VSS.n1936 VSS.n1182 25.6005
R3234 VSS.n1942 VSS.n1183 25.6005
R3235 VSS.n1954 VSS.n1953 25.6005
R3236 VSS.n935 VSS.n931 25.6005
R3237 VSS.n2108 VSS.n876 25.6005
R3238 VSS.n2108 VSS.n2107 25.6005
R3239 VSS.n2107 VSS.n2106 25.6005
R3240 VSS.n2106 VSS.n877 25.6005
R3241 VSS.n893 VSS.n877 25.6005
R3242 VSS.n2092 VSS.n893 25.6005
R3243 VSS.n2092 VSS.n2091 25.6005
R3244 VSS.n2091 VSS.n2090 25.6005
R3245 VSS.n2090 VSS.n894 25.6005
R3246 VSS.n2084 VSS.n894 25.6005
R3247 VSS.n2084 VSS.n2083 25.6005
R3248 VSS.n2011 VSS.n2010 25.6005
R3249 VSS.n2010 VSS.n2009 25.6005
R3250 VSS.n2009 VSS.n2006 25.6005
R3251 VSS.n2006 VSS.n2005 25.6005
R3252 VSS.n2005 VSS.n2002 25.6005
R3253 VSS.n2002 VSS.n2001 25.6005
R3254 VSS.n2001 VSS.n1998 25.6005
R3255 VSS.n1998 VSS.n1997 25.6005
R3256 VSS.n1997 VSS.n1994 25.6005
R3257 VSS.n1994 VSS.n1993 25.6005
R3258 VSS.n1993 VSS.n1990 25.6005
R3259 VSS.n1990 VSS.n1989 25.6005
R3260 VSS.n1989 VSS.n1986 25.6005
R3261 VSS.n1986 VSS.n1985 25.6005
R3262 VSS.n1985 VSS.n1982 25.6005
R3263 VSS.n1982 VSS.n1981 25.6005
R3264 VSS.n1981 VSS.n1978 25.6005
R3265 VSS.n1978 VSS.n1977 25.6005
R3266 VSS.n1977 VSS.n1974 25.6005
R3267 VSS.n1974 VSS.n1973 25.6005
R3268 VSS.n1973 VSS.n1971 25.6005
R3269 VSS.n1971 VSS.n924 25.6005
R3270 VSS.n2018 VSS.n2017 25.6005
R3271 VSS.n2021 VSS.n2018 25.6005
R3272 VSS.n2022 VSS.n2021 25.6005
R3273 VSS.n2023 VSS.n2022 25.6005
R3274 VSS.n2028 VSS.n2023 25.6005
R3275 VSS.n2029 VSS.n2028 25.6005
R3276 VSS.n2031 VSS.n2029 25.6005
R3277 VSS.n2032 VSS.n2031 25.6005
R3278 VSS.n2033 VSS.n2032 25.6005
R3279 VSS.n2034 VSS.n2033 25.6005
R3280 VSS.n2035 VSS.n2034 25.6005
R3281 VSS.n2082 VSS.n901 25.6005
R3282 VSS.n2077 VSS.n901 25.6005
R3283 VSS.n2077 VSS.n2076 25.6005
R3284 VSS.n2076 VSS.n2075 25.6005
R3285 VSS.n2075 VSS.n2072 25.6005
R3286 VSS.n2072 VSS.n2071 25.6005
R3287 VSS.n920 VSS.n915 25.6005
R3288 VSS.n2060 VSS.n2059 25.6005
R3289 VSS.n2054 VSS.n2051 25.6005
R3290 VSS.n2051 VSS.n2050 25.6005
R3291 VSS.n2050 VSS.n2047 25.6005
R3292 VSS.n2047 VSS.n2046 25.6005
R3293 VSS.n2046 VSS.n2043 25.6005
R3294 VSS.n2043 VSS.n2042 25.6005
R3295 VSS.n2042 VSS.n2039 25.6005
R3296 VSS.n2039 VSS.n2038 25.6005
R3297 VSS.n550 VSS.n545 25.6005
R3298 VSS.n550 VSS.n549 25.6005
R3299 VSS.n556 VSS.n549 25.6005
R3300 VSS.n557 VSS.n556 25.6005
R3301 VSS.n563 VSS.n562 25.6005
R3302 VSS.n564 VSS.n563 25.6005
R3303 VSS.n564 VSS.n537 25.6005
R3304 VSS.n575 VSS.n537 25.6005
R3305 VSS.n576 VSS.n575 25.6005
R3306 VSS.n577 VSS.n576 25.6005
R3307 VSS.n577 VSS.n448 25.6005
R3308 VSS.n2291 VSS.n448 25.6005
R3309 VSS.n2291 VSS.n2290 25.6005
R3310 VSS.n2290 VSS.n2289 25.6005
R3311 VSS.n2289 VSS.n449 25.6005
R3312 VSS.n2283 VSS.n449 25.6005
R3313 VSS.n2283 VSS.n2282 25.6005
R3314 VSS.n2282 VSS.n2281 25.6005
R3315 VSS.n2281 VSS.n456 25.6005
R3316 VSS.n2275 VSS.n456 25.6005
R3317 VSS.n2275 VSS.n2274 25.6005
R3318 VSS.n2274 VSS.n2273 25.6005
R3319 VSS.n2273 VSS.n463 25.6005
R3320 VSS.n2267 VSS.n463 25.6005
R3321 VSS.n2267 VSS.n2266 25.6005
R3322 VSS.n2266 VSS.n2265 25.6005
R3323 VSS.n2265 VSS.n470 25.6005
R3324 VSS.n2259 VSS.n470 25.6005
R3325 VSS.n2259 VSS.n2258 25.6005
R3326 VSS.n2258 VSS.n2257 25.6005
R3327 VSS.n2257 VSS.n477 25.6005
R3328 VSS.n2251 VSS.n477 25.6005
R3329 VSS.n2251 VSS.n2250 25.6005
R3330 VSS.n2250 VSS.n2249 25.6005
R3331 VSS.n2249 VSS.n484 25.6005
R3332 VSS.n2243 VSS.n484 25.6005
R3333 VSS.n2243 VSS.n2242 25.6005
R3334 VSS.n2242 VSS.n2241 25.6005
R3335 VSS.n2241 VSS.n491 25.6005
R3336 VSS.n2235 VSS.n491 25.6005
R3337 VSS.n2235 VSS.n2234 25.6005
R3338 VSS.n2234 VSS.n2233 25.6005
R3339 VSS.n2233 VSS.n498 25.6005
R3340 VSS.n2227 VSS.n498 25.6005
R3341 VSS.n2227 VSS.n2226 25.6005
R3342 VSS.n2226 VSS.n2225 25.6005
R3343 VSS.n2225 VSS.n505 25.6005
R3344 VSS.n2219 VSS.n505 25.6005
R3345 VSS.n2219 VSS.n2218 25.6005
R3346 VSS.n2218 VSS.n2217 25.6005
R3347 VSS.n2217 VSS.n512 25.6005
R3348 VSS.n2211 VSS.n512 25.6005
R3349 VSS.n2211 VSS.n2210 25.6005
R3350 VSS.n2210 VSS.n2209 25.6005
R3351 VSS.n2209 VSS.n519 25.6005
R3352 VSS.n2203 VSS.n519 25.6005
R3353 VSS.n2203 VSS.n2202 25.6005
R3354 VSS.n2197 VSS.n528 25.6005
R3355 VSS.n532 VSS.n528 25.6005
R3356 VSS.n641 VSS.n532 25.6005
R3357 VSS.n558 VSS.n541 25.6005
R3358 VSS.n568 VSS.n541 25.6005
R3359 VSS.n569 VSS.n568 25.6005
R3360 VSS.n571 VSS.n569 25.6005
R3361 VSS.n571 VSS.n570 25.6005
R3362 VSS.n570 VSS.n533 25.6005
R3363 VSS.n582 VSS.n533 25.6005
R3364 VSS.n583 VSS.n582 25.6005
R3365 VSS.n585 VSS.n583 25.6005
R3366 VSS.n586 VSS.n585 25.6005
R3367 VSS.n587 VSS.n586 25.6005
R3368 VSS.n588 VSS.n587 25.6005
R3369 VSS.n590 VSS.n588 25.6005
R3370 VSS.n591 VSS.n590 25.6005
R3371 VSS.n592 VSS.n591 25.6005
R3372 VSS.n593 VSS.n592 25.6005
R3373 VSS.n595 VSS.n593 25.6005
R3374 VSS.n596 VSS.n595 25.6005
R3375 VSS.n597 VSS.n596 25.6005
R3376 VSS.n598 VSS.n597 25.6005
R3377 VSS.n600 VSS.n598 25.6005
R3378 VSS.n601 VSS.n600 25.6005
R3379 VSS.n602 VSS.n601 25.6005
R3380 VSS.n603 VSS.n602 25.6005
R3381 VSS.n605 VSS.n603 25.6005
R3382 VSS.n606 VSS.n605 25.6005
R3383 VSS.n608 VSS.n606 25.6005
R3384 VSS.n609 VSS.n608 25.6005
R3385 VSS.n611 VSS.n609 25.6005
R3386 VSS.n612 VSS.n611 25.6005
R3387 VSS.n613 VSS.n612 25.6005
R3388 VSS.n614 VSS.n613 25.6005
R3389 VSS.n616 VSS.n614 25.6005
R3390 VSS.n617 VSS.n616 25.6005
R3391 VSS.n618 VSS.n617 25.6005
R3392 VSS.n619 VSS.n618 25.6005
R3393 VSS.n621 VSS.n619 25.6005
R3394 VSS.n622 VSS.n621 25.6005
R3395 VSS.n623 VSS.n622 25.6005
R3396 VSS.n624 VSS.n623 25.6005
R3397 VSS.n626 VSS.n624 25.6005
R3398 VSS.n627 VSS.n626 25.6005
R3399 VSS.n628 VSS.n627 25.6005
R3400 VSS.n629 VSS.n628 25.6005
R3401 VSS.n631 VSS.n629 25.6005
R3402 VSS.n632 VSS.n631 25.6005
R3403 VSS.n633 VSS.n632 25.6005
R3404 VSS.n634 VSS.n633 25.6005
R3405 VSS.n636 VSS.n634 25.6005
R3406 VSS.n637 VSS.n636 25.6005
R3407 VSS.n638 VSS.n637 25.6005
R3408 VSS.n639 VSS.n638 25.6005
R3409 VSS.n640 VSS.n639 25.6005
R3410 VSS.n745 VSS.n743 25.6005
R3411 VSS.n743 VSS.n740 25.6005
R3412 VSS.n740 VSS.n739 25.6005
R3413 VSS.n739 VSS.n736 25.6005
R3414 VSS.n736 VSS.n735 25.6005
R3415 VSS.n735 VSS.n732 25.6005
R3416 VSS.n732 VSS.n731 25.6005
R3417 VSS.n731 VSS.n728 25.6005
R3418 VSS.n728 VSS.n727 25.6005
R3419 VSS.n727 VSS.n724 25.6005
R3420 VSS.n724 VSS.n723 25.6005
R3421 VSS.n723 VSS.n720 25.6005
R3422 VSS.n720 VSS.n719 25.6005
R3423 VSS.n719 VSS.n716 25.6005
R3424 VSS.n716 VSS.n715 25.6005
R3425 VSS.n715 VSS.n712 25.6005
R3426 VSS.n712 VSS.n711 25.6005
R3427 VSS.n711 VSS.n708 25.6005
R3428 VSS.n708 VSS.n707 25.6005
R3429 VSS.n707 VSS.n704 25.6005
R3430 VSS.n704 VSS.n697 25.6005
R3431 VSS.n2160 VSS.n697 25.6005
R3432 VSS.n2154 VSS.n746 25.6005
R3433 VSS.n2154 VSS.n2153 25.6005
R3434 VSS.n2153 VSS.n2152 25.6005
R3435 VSS.n2152 VSS.n747 25.6005
R3436 VSS.n762 VSS.n747 25.6005
R3437 VSS.n2140 VSS.n762 25.6005
R3438 VSS.n2140 VSS.n2139 25.6005
R3439 VSS.n2139 VSS.n2138 25.6005
R3440 VSS.n2138 VSS.n763 25.6005
R3441 VSS.n778 VSS.n763 25.6005
R3442 VSS.n2126 VSS.n778 25.6005
R3443 VSS.n2125 VSS.n2124 25.6005
R3444 VSS.n2124 VSS.n779 25.6005
R3445 VSS.n793 VSS.n779 25.6005
R3446 VSS.n794 VSS.n793 25.6005
R3447 VSS.n797 VSS.n794 25.6005
R3448 VSS.n798 VSS.n797 25.6005
R3449 VSS.n801 VSS.n798 25.6005
R3450 VSS.n802 VSS.n801 25.6005
R3451 VSS.n805 VSS.n802 25.6005
R3452 VSS.n806 VSS.n805 25.6005
R3453 VSS.n809 VSS.n806 25.6005
R3454 VSS.n810 VSS.n809 25.6005
R3455 VSS.n813 VSS.n810 25.6005
R3456 VSS.n814 VSS.n813 25.6005
R3457 VSS.n817 VSS.n814 25.6005
R3458 VSS.n818 VSS.n817 25.6005
R3459 VSS.n821 VSS.n818 25.6005
R3460 VSS.n822 VSS.n821 25.6005
R3461 VSS.n825 VSS.n822 25.6005
R3462 VSS.n827 VSS.n825 25.6005
R3463 VSS.n828 VSS.n827 25.6005
R3464 VSS.n856 VSS.n828 25.6005
R3465 VSS.n2159 VSS.n2158 25.6005
R3466 VSS.n838 VSS.n837 25.6005
R3467 VSS.n844 VSS.n831 25.6005
R3468 VSS.n854 VSS.n851 25.6005
R3469 VSS.n855 VSS.n854 25.6005
R3470 VSS.t25 VSS.n2086 25.0064
R3471 VSS.n2295 VSS.n2293 24.8841
R3472 VSS.n310 VSS.n304 24.8476
R3473 VSS.n365 VSS.n359 24.8476
R3474 VSS.n65 VSS.n47 24.8476
R3475 VSS.n19 VSS.n18 24.8476
R3476 VSS.n293 VSS.n230 24.8476
R3477 VSS.n2510 VSS.n2509 24.8476
R3478 VSS.n1761 VSS.n1423 24.8476
R3479 VSS.n1278 VSS.n1277 24.8476
R3480 VSS.n1210 VSS.n1207 24.8476
R3481 VSS.n1369 VSS.n1339 24.8476
R3482 VSS.n1850 VSS.n1848 24.8476
R3483 VSS.n1901 VSS.n1325 24.8476
R3484 VSS.n1891 VSS.n756 24.8476
R3485 VSS.n1909 VSS.n1299 24.8476
R3486 VSS.n1918 VSS.n1193 24.8476
R3487 VSS.n60 VSS.n59 24.75
R3488 VSS.n23 VSS.n22 24.75
R3489 VSS.n323 VSS.n299 24.2609
R3490 VSS.n317 VSS.n297 24.2609
R3491 VSS.n378 VSS.n372 24.2609
R3492 VSS.n383 VSS.n374 24.2609
R3493 VSS.n53 VSS.n49 24.2609
R3494 VSS.n27 VSS.n6 24.2609
R3495 VSS.n274 VSS.n272 23.7181
R3496 VSS.n281 VSS.n236 23.7181
R3497 VSS.n2525 VSS.n2499 23.7181
R3498 VSS.n2521 VSS.n2500 23.7181
R3499 VSS.n2201 VSS.n526 23.7181
R3500 VSS.n2164 VSS.n680 23.4436
R3501 VSS.n323 VSS.n300 23.3417
R3502 VSS.n317 VSS.n298 23.3417
R3503 VSS.n307 VSS.n303 23.3417
R3504 VSS.n378 VSS.n373 23.3417
R3505 VSS.n383 VSS.n375 23.3417
R3506 VSS.n362 VSS.n358 23.3417
R3507 VSS.n69 VSS.n68 23.3417
R3508 VSS.n53 VSS.n50 23.3417
R3509 VSS.n28 VSS.n27 23.3417
R3510 VSS.n15 VSS.n10 23.3417
R3511 VSS.n1274 VSS.n1248 23.3417
R3512 VSS.n1211 VSS.n1205 23.3417
R3513 VSS.n1368 VSS.n1341 23.3417
R3514 VSS.n1854 VSS.n1853 23.3417
R3515 VSS.n1821 VSS.n1817 22.9652
R3516 VSS.n2117 VSS.n2116 22.9652
R3517 VSS.n2175 VSS.n2174 22.9652
R3518 VSS.n1943 VSS.n1182 22.9652
R3519 VSS.n2068 VSS.n914 22.9652
R3520 VSS.n2111 VSS.n2110 22.9226
R3521 VSS.n2104 VSS.n879 22.9226
R3522 VSS.n2024 VSS.n888 22.9226
R3523 VSS.n311 VSS.n310 22.4252
R3524 VSS.n366 VSS.n365 22.4252
R3525 VSS.n2308 VSS.t26 22.4016
R3526 VSS.n2444 VSS.t43 22.4016
R3527 VSS.n327 VSS.n326 21.8358
R3528 VSS.n330 VSS.n296 21.8358
R3529 VSS.n313 VSS.n302 21.8358
R3530 VSS.n390 VSS.n371 21.8358
R3531 VSS.n387 VSS.n386 21.8358
R3532 VSS.n368 VSS.n357 21.8358
R3533 VSS.n71 VSS.n45 21.8358
R3534 VSS.n57 VSS.n56 21.8358
R3535 VSS.n30 VSS.n5 21.8358
R3536 VSS.n14 VSS.n11 21.8358
R3537 VSS.n1757 VSS.n1424 21.8358
R3538 VSS.n1273 VSS.n1250 21.8358
R3539 VSS.n1215 VSS.n1214 21.8358
R3540 VSS.n1365 VSS.n1364 21.8358
R3541 VSS.n1857 VSS.n1846 21.8358
R3542 VSS.n1819 VSS.n1394 21.8358
R3543 VSS.n2114 VSS.n2113 21.8358
R3544 VSS.n2178 VSS.n2177 21.8358
R3545 VSS.n1954 VSS.n930 21.8358
R3546 VSS.n834 VSS.n698 21.8358
R3547 VSS.n2372 VSS.t33 21.3597
R3548 VSS.t9 VSS.n157 21.3597
R3549 VSS.n286 VSS.n284 21.0829
R3550 VSS.n396 VSS.n230 21.0829
R3551 VSS.n2514 VSS.n2502 21.0829
R3552 VSS.n2509 VSS.n2507 21.0829
R3553 VSS.n1835 VSS.n1393 21.0829
R3554 VSS.n1885 VSS.n883 21.0829
R3555 VSS.n664 VSS.n660 21.0829
R3556 VSS.n1952 VSS.n931 21.0829
R3557 VSS.n1906 VSS.n701 20.4928
R3558 VSS.n1270 VSS.n1269 20.3299
R3559 VSS.n1218 VSS.n1203 20.3299
R3560 VSS.n1361 VSS.n1343 20.3299
R3561 VSS.n1858 VSS.n1844 20.3299
R3562 VSS.n1733 VSS.n1732 20.3299
R3563 VSS.n2100 VSS.n884 20.3299
R3564 VSS.n2186 VSS.n658 20.3299
R3565 VSS.n1178 VSS.n1177 20.3299
R3566 VSS.n2328 VSS.t3 20.3178
R3567 VSS.n133 VSS.t47 20.3178
R3568 VSS.n2025 VSS.t40 20.3178
R3569 VSS.n286 VSS.n285 19.9534
R3570 VSS.n2514 VSS.n2513 19.9534
R3571 VSS.n1329 VSS.n1328 19.7969
R3572 VSS.n2156 VSS.n700 19.7969
R3573 VSS.n2150 VSS.n749 19.7969
R3574 VSS.n2149 VSS.n751 19.7969
R3575 VSS.n841 VSS.n840 19.7969
R3576 VSS.n829 VSS.n759 19.7969
R3577 VSS.n2136 VSS.n765 19.7969
R3578 VSS.n2135 VSS.n767 19.7969
R3579 VSS.n1187 VSS.n773 19.7969
R3580 VSS.n2129 VSS.n2128 19.7969
R3581 VSS.n1754 VSS.n1753 18.824
R3582 VSS.n1266 VSS.n1252 18.824
R3583 VSS.n1219 VSS.n1201 18.824
R3584 VSS.n1360 VSS.n1345 18.824
R3585 VSS.n1862 VSS.n1861 18.824
R3586 VSS.n1657 VSS.n1656 18.7549
R3587 VSS.n1736 VSS.n1735 18.7549
R3588 VSS.n1743 VSS.n1742 18.7549
R3589 VSS.n1831 VSS.n1398 18.7549
R3590 VSS.n1825 VSS.n1824 18.7549
R3591 VSS.n1813 VSS.n1409 18.7549
R3592 VSS.n1763 VSS.n1423 18.5363
R3593 VSS.n1332 VSS.n1331 18.4476
R3594 VSS.n1892 VSS.n770 18.4476
R3595 VSS.n1313 VSS.n1298 18.4476
R3596 VSS.n1926 VSS.n1189 18.4476
R3597 VSS.n2067 VSS.n915 18.4476
R3598 VSS.t17 VSS.n2120 18.234
R3599 VSS.n2064 VSS.n2063 18.0711
R3600 VSS.n850 VSS.n849 18.0711
R3601 VSS.n1744 VSS.t6 17.713
R3602 VSS.t21 VSS.n2142 17.713
R3603 VSS.t19 VSS.n2094 17.713
R3604 VSS.n273 VSS.n236 17.3181
R3605 VSS.n2524 VSS.n2500 17.3181
R3606 VSS.n1265 VSS.n1254 17.3181
R3607 VSS.n1224 VSS.n1223 17.3181
R3608 VSS.n1357 VSS.n1356 17.3181
R3609 VSS.n1865 VSS.n1842 17.3181
R3610 VSS.n837 VSS.n836 17.3181
R3611 VSS.n1258 VSS.n1257 17.1928
R3612 VSS.n1230 VSS.n1229 17.1928
R3613 VSS.n1350 VSS.n1349 17.1928
R3614 VSS.n1870 VSS.n1838 17.1928
R3615 VSS.t16 VSS.n2170 17.1921
R3616 VSS.n2056 VSS.n2055 16.9417
R3617 VSS.n843 VSS.n833 16.9417
R3618 VSS.n1735 VSS.n1432 16.6711
R3619 VSS.n1742 VSS.n1427 16.6711
R3620 VSS.n1744 VSS.n1743 16.6711
R3621 VSS.n1832 VSS.n1831 16.6711
R3622 VSS.n1751 VSS.n1398 16.6711
R3623 VSS.n1825 VSS.n1404 16.6711
R3624 VSS.n1824 VSS.n1406 16.6711
R3625 VSS.n1814 VSS.n1813 16.6711
R3626 VSS.n1409 VSS.n673 16.6711
R3627 VSS.n1432 VSS.t0 16.1502
R3628 VSS.n1262 VSS.n1261 15.8123
R3629 VSS.n1227 VSS.n1199 15.8123
R3630 VSS.n1353 VSS.n1347 15.8123
R3631 VSS.n1866 VSS.n1840 15.8123
R3632 VSS.n1328 VSS.n700 15.6292
R3633 VSS.n1905 VSS.n749 15.6292
R3634 VSS.n2150 VSS.n2149 15.6292
R3635 VSS.n840 VSS.n751 15.6292
R3636 VSS.n2142 VSS.n759 15.6292
R3637 VSS.n829 VSS.n765 15.6292
R3638 VSS.n2136 VSS.n2135 15.6292
R3639 VSS.n2129 VSS.n773 15.6292
R3640 VSS.n2128 VSS.n775 15.6292
R3641 VSS.n2321 VSS.t3 15.1082
R3642 VSS.n2432 VSS.t47 15.1082
R3643 VSS.n2121 VSS.n781 15.1082
R3644 VSS.n327 VSS.n316 14.5711
R3645 VSS.n331 VSS.n330 14.5711
R3646 VSS.n314 VSS.n313 14.5711
R3647 VSS.n391 VSS.n390 14.5711
R3648 VSS.n387 VSS.n376 14.5711
R3649 VSS.n369 VSS.n368 14.5711
R3650 VSS.n72 VSS.n71 14.5711
R3651 VSS.n57 VSS.n51 14.5711
R3652 VSS.n31 VSS.n30 14.5711
R3653 VSS.n11 VSS.n3 14.5711
R3654 VSS.n1748 VSS.n1747 14.3064
R3655 VSS.n1258 VSS.n1256 14.3064
R3656 VSS.n1229 VSS.n1228 14.3064
R3657 VSS.n1352 VSS.n1349 14.3064
R3658 VSS.n1870 VSS.n1869 14.3064
R3659 VSS.t33 VSS.n165 14.0663
R3660 VSS.n2384 VSS.t9 14.0663
R3661 VSS.n1729 VSS.n1728 13.9299
R3662 VSS.n2098 VSS.n2097 13.9299
R3663 VSS.n2189 VSS.n2188 13.9299
R3664 VSS.n952 VSS.n934 13.9299
R3665 VSS.n2060 VSS.n921 13.5534
R3666 VSS.n848 VSS.n831 13.5534
R3667 VSS.t15 VSS.n2162 13.5454
R3668 VSS.n2056 VSS.n923 13.177
R3669 VSS.n2198 VSS.n526 13.177
R3670 VSS.n845 VSS.n843 13.177
R3671 VSS.n2315 VSS.t26 13.0244
R3672 VSS.n125 VSS.t43 13.0244
R3673 VSS.t18 VSS.n871 13.0244
R3674 VSS.n2111 VSS.n871 12.5035
R3675 VSS.n2110 VSS.n873 12.5035
R3676 VSS.t51 VSS.n873 12.5035
R3677 VSS.n2019 VSS.n879 12.5035
R3678 VSS.n2104 VSS.n2103 12.5035
R3679 VSS.n2025 VSS.n2024 12.5035
R3680 VSS.n2095 VSS.n888 12.5035
R3681 VSS.n2059 VSS.n923 12.424
R3682 VSS.n2198 VSS.n2197 12.424
R3683 VSS.n845 VSS.n844 12.424
R3684 VSS.n2063 VSS.n921 12.0476
R3685 VSS.n849 VSS.n848 12.0476
R3686 VSS.n680 VSS.n674 11.9825
R3687 VSS.n841 VSS.t23 11.9825
R3688 VSS.n1733 VSS.n1729 11.6711
R3689 VSS.n2098 VSS.n884 11.6711
R3690 VSS.n2188 VSS.n658 11.6711
R3691 VSS.n1177 VSS.n934 11.6711
R3692 VSS.n1753 VSS.n1748 11.2946
R3693 VSS.n1261 VSS.n1256 11.2946
R3694 VSS.n1228 VSS.n1227 11.2946
R3695 VSS.n1353 VSS.n1352 11.2946
R3696 VSS.n1869 VSS.n1840 11.2946
R3697 VSS.n1381 VSS.n1375 11.0636
R3698 VSS.n1380 VSS.n1376 11.0636
R3699 VSS.n1379 VSS.n1377 11.0636
R3700 VSS.n1378 VSS.n1373 11.0636
R3701 VSS.n1877 VSS.n1382 11.0636
R3702 VSS.n1876 VSS.n1383 11.0636
R3703 VSS.n1875 VSS.n1384 11.0636
R3704 VSS.n1874 VSS.n1385 11.0636
R3705 VSS.n1873 VSS.n1872 11.0636
R3706 VSS.n1282 VSS.n1281 11.0636
R3707 VSS.n1283 VSS.n1245 11.0636
R3708 VSS.n1284 VSS.n1244 11.0636
R3709 VSS.n1285 VSS.n1235 11.0636
R3710 VSS.n1291 VSS.n1231 11.0636
R3711 VSS.n1290 VSS.n1232 11.0636
R3712 VSS.n1289 VSS.n1233 11.0636
R3713 VSS.n1288 VSS.n1234 11.0636
R3714 VSS.n1287 VSS.n1286 11.0636
R3715 VSS.n2163 VSS.t15 10.9406
R3716 VSS.n2162 VSS.n694 10.9406
R3717 VSS.n1736 VSS.t24 10.4196
R3718 VSS.t20 VSS.n1406 10.4196
R3719 VSS.t57 VSS.n1905 10.4196
R3720 VSS.n2019 VSS.t51 10.4196
R3721 VSS.n2087 VSS.t25 10.4196
R3722 VSS.n1906 VSS.t5 10.2467
R3723 VSS.n1921 VSS.t23 10.2467
R3724 VSS.t22 VSS.n1404 9.89868
R3725 VSS.n1957 VSS.t18 9.89868
R3726 VSS.n1262 VSS.n1254 9.78874
R3727 VSS.n1224 VSS.n1199 9.78874
R3728 VSS.n1356 VSS.n1347 9.78874
R3729 VSS.n1866 VSS.n1865 9.78874
R3730 VSS.n1278 VSS.n1246 9.58499
R3731 VSS.n1208 VSS.n1207 9.58499
R3732 VSS.n1371 VSS.n1339 9.58499
R3733 VSS.n1850 VSS.n1849 9.58499
R3734 VSS.n2199 VSS.n528 9.52595
R3735 VSS.n2523 VSS.n2499 9.49023
R3736 VSS.n272 VSS.n235 9.49023
R3737 VSS.n1179 VSS.n934 9.49023
R3738 VSS.n1944 VSS.n1943 9.49023
R3739 VSS.n1917 VSS.n1189 9.49023
R3740 VSS.n1910 VSS.n1298 9.49023
R3741 VSS.n1900 VSS.n1332 9.49023
R3742 VSS.n1893 VSS.n1892 9.49023
R3743 VSS.n2116 VSS.n2115 9.49023
R3744 VSS.n2099 VSS.n2098 9.49023
R3745 VSS.n1821 VSS.n1820 9.49023
R3746 VSS.n1731 VSS.n1729 9.49023
R3747 VSS.n2176 VSS.n2175 9.49023
R3748 VSS.n2188 VSS.n2187 9.49023
R3749 VSS.n1755 VSS.n1748 9.41955
R3750 VSS.n835 VSS.n698 9.41955
R3751 VSS.n850 VSS.n1 9.35854
R3752 VSS.n318 VSS.n317 9.3005
R3753 VSS.n296 VSS.n295 9.3005
R3754 VSS.n310 VSS.n309 9.3005
R3755 VSS.n308 VSS.n307 9.3005
R3756 VSS.n302 VSS.n301 9.3005
R3757 VSS.n324 VSS.n323 9.3005
R3758 VSS.n326 VSS.n325 9.3005
R3759 VSS.n384 VSS.n383 9.3005
R3760 VSS.n386 VSS.n385 9.3005
R3761 VSS.n365 VSS.n364 9.3005
R3762 VSS.n363 VSS.n362 9.3005
R3763 VSS.n357 VSS.n356 9.3005
R3764 VSS.n379 VSS.n378 9.3005
R3765 VSS.n371 VSS.n370 9.3005
R3766 VSS.n54 VSS.n53 9.3005
R3767 VSS.n56 VSS.n55 9.3005
R3768 VSS.n66 VSS.n65 9.3005
R3769 VSS.n68 VSS.n67 9.3005
R3770 VSS.n45 VSS.n44 9.3005
R3771 VSS.n19 VSS.n9 9.3005
R3772 VSS.n12 VSS.n10 9.3005
R3773 VSS.n14 VSS.n13 9.3005
R3774 VSS.n27 VSS.n26 9.3005
R3775 VSS.n5 VSS.n4 9.3005
R3776 VSS.n396 VSS.n395 9.3005
R3777 VSS.n285 VSS.n231 9.3005
R3778 VSS.n282 VSS.n281 9.3005
R3779 VSS.n394 VSS.n228 9.3005
R3780 VSS.n294 VSS.n293 9.3005
R3781 VSS.n284 VSS.n283 9.3005
R3782 VSS.n273 VSS.n235 9.3005
R3783 VSS.n2507 VSS.n75 9.3005
R3784 VSS.n2513 VSS.n2512 9.3005
R3785 VSS.n2522 VSS.n2521 9.3005
R3786 VSS.n2524 VSS.n2523 9.3005
R3787 VSS.n2502 VSS.n2501 9.3005
R3788 VSS.n2511 VSS.n2510 9.3005
R3789 VSS.n2560 VSS.n2559 9.3005
R3790 VSS.n1755 VSS.n1754 9.3005
R3791 VSS.n1757 VSS.n1756 9.3005
R3792 VSS.n1762 VSS.n1761 9.3005
R3793 VSS.n1279 VSS.n1278 9.3005
R3794 VSS.n1248 VSS.n1247 9.3005
R3795 VSS.n1273 VSS.n1272 9.3005
R3796 VSS.n1271 VSS.n1270 9.3005
R3797 VSS.n1252 VSS.n1251 9.3005
R3798 VSS.n1265 VSS.n1264 9.3005
R3799 VSS.n1263 VSS.n1262 9.3005
R3800 VSS.n1256 VSS.n1255 9.3005
R3801 VSS.n1207 VSS.n1206 9.3005
R3802 VSS.n1212 VSS.n1211 9.3005
R3803 VSS.n1214 VSS.n1213 9.3005
R3804 VSS.n1203 VSS.n1202 9.3005
R3805 VSS.n1220 VSS.n1219 9.3005
R3806 VSS.n1223 VSS.n1222 9.3005
R3807 VSS.n1221 VSS.n1199 9.3005
R3808 VSS.n1228 VSS.n1198 9.3005
R3809 VSS.n1339 VSS.n1338 9.3005
R3810 VSS.n1368 VSS.n1367 9.3005
R3811 VSS.n1366 VSS.n1365 9.3005
R3812 VSS.n1343 VSS.n1342 9.3005
R3813 VSS.n1360 VSS.n1359 9.3005
R3814 VSS.n1358 VSS.n1357 9.3005
R3815 VSS.n1347 VSS.n1346 9.3005
R3816 VSS.n1352 VSS.n1351 9.3005
R3817 VSS.n1851 VSS.n1850 9.3005
R3818 VSS.n1853 VSS.n1852 9.3005
R3819 VSS.n1846 VSS.n1845 9.3005
R3820 VSS.n1859 VSS.n1858 9.3005
R3821 VSS.n1861 VSS.n1860 9.3005
R3822 VSS.n1842 VSS.n1841 9.3005
R3823 VSS.n1867 VSS.n1866 9.3005
R3824 VSS.n1869 VSS.n1868 9.3005
R3825 VSS.n1732 VSS.n1731 9.3005
R3826 VSS.n1836 VSS.n1835 9.3005
R3827 VSS.n1820 VSS.n1819 9.3005
R3828 VSS.n1901 VSS.n1900 9.3005
R3829 VSS.n2100 VSS.n2099 9.3005
R3830 VSS.n1886 VSS.n1885 9.3005
R3831 VSS.n2115 VSS.n2114 9.3005
R3832 VSS.n1893 VSS.n756 9.3005
R3833 VSS.n2147 VSS.n755 9.3005
R3834 VSS.n1910 VSS.n1909 9.3005
R3835 VSS.n1320 VSS.n1194 9.3005
R3836 VSS.n1918 VSS.n1917 9.3005
R3837 VSS.n1944 VSS.n930 9.3005
R3838 VSS.n1952 VSS.n1951 9.3005
R3839 VSS.n1179 VSS.n1178 9.3005
R3840 VSS.n2177 VSS.n2176 9.3005
R3841 VSS.n1293 VSS.n664 9.3005
R3842 VSS.n2187 VSS.n2186 9.3005
R3843 VSS.n2055 VSS.n0 9.3005
R3844 VSS.n916 VSS.n914 9.3005
R3845 VSS.n2067 VSS.n2066 9.3005
R3846 VSS.n2065 VSS.n2064 9.3005
R3847 VSS.n921 VSS.n917 9.3005
R3848 VSS.n923 VSS.n922 9.3005
R3849 VSS.n2199 VSS.n2198 9.3005
R3850 VSS.n2201 VSS.n2200 9.3005
R3851 VSS.n846 VSS.n845 9.3005
R3852 VSS.n848 VSS.n847 9.3005
R3853 VSS.n833 VSS.n832 9.3005
R3854 VSS.n836 VSS.n835 9.3005
R3855 VSS.n1751 VSS.t22 8.85676
R3856 VSS.n2055 VSS.n2054 8.65932
R3857 VSS.n838 VSS.n833 8.65932
R3858 VSS.n1814 VSS.t20 8.33581
R3859 VSS.n2156 VSS.n701 8.33581
R3860 VSS.n274 VSS.n273 8.28285
R3861 VSS.n2525 VSS.n2524 8.28285
R3862 VSS.n1266 VSS.n1265 8.28285
R3863 VSS.n1223 VSS.n1201 8.28285
R3864 VSS.n1357 VSS.n1345 8.28285
R3865 VSS.n1862 VSS.n1842 8.28285
R3866 VSS.n836 VSS.n834 8.28285
R3867 VSS.n311 VSS.n306 8.2073
R3868 VSS.n366 VSS.n361 8.2073
R3869 VSS.n2334 VSS.t30 7.81485
R3870 VSS.n2420 VSS.t1 7.81485
R3871 VSS.n2013 VSS.n1959 7.81485
R3872 VSS.n2064 VSS.n920 7.52991
R3873 VSS.n851 VSS.n850 7.52991
R3874 VSS.n2183 VSS.t0 7.3192
R3875 VSS.n938 VSS.t40 7.3192
R3876 VSS.n1904 VSS.n701 7.29389
R3877 VSS.n2254 VSS.n480 7.24494
R3878 VSS.n1332 VSS.n1325 7.15344
R3879 VSS.n1892 VSS.n1891 7.15344
R3880 VSS.n1299 VSS.n1298 7.15344
R3881 VSS.n1193 VSS.n1189 7.15344
R3882 VSS.n2068 VSS.n2067 7.15344
R3883 VSS.n1754 VSS.n1424 6.77697
R3884 VSS.n1269 VSS.n1252 6.77697
R3885 VSS.n1219 VSS.n1218 6.77697
R3886 VSS.n1361 VSS.n1360 6.77697
R3887 VSS.n1861 VSS.n1844 6.77697
R3888 VSS.t13 VSS.n173 6.77294
R3889 VSS.n2396 VSS.t45 6.77294
R3890 VSS.n322 VSS.n299 6.41949
R3891 VSS.n319 VSS.n297 6.41949
R3892 VSS.n380 VSS.n372 6.41949
R3893 VSS.n382 VSS.n374 6.41949
R3894 VSS.n52 VSS.n49 6.41949
R3895 VSS.n25 VSS.n6 6.41949
R3896 VSS.n1656 VSS.t24 6.25198
R3897 VSS.t122 VSS.n328 5.8005
R3898 VSS.n328 VSS.t80 5.8005
R3899 VSS.n329 VSS.t44 5.8005
R3900 VSS.n329 VSS.t122 5.8005
R3901 VSS.n312 VSS.t37 5.8005
R3902 VSS.n312 VSS.t73 5.8005
R3903 VSS.n389 VSS.t90 5.8005
R3904 VSS.n389 VSS.t88 5.8005
R3905 VSS.t88 VSS.n388 5.8005
R3906 VSS.n388 VSS.t49 5.8005
R3907 VSS.n367 VSS.t84 5.8005
R3908 VSS.n367 VSS.t53 5.8005
R3909 VSS.n333 VSS.t129 5.8005
R3910 VSS.n333 VSS.t136 5.8005
R3911 VSS.n337 VSS.t12 5.8005
R3912 VSS.n337 VSS.t54 5.8005
R3913 VSS.n341 VSS.t39 5.8005
R3914 VSS.n341 VSS.t135 5.8005
R3915 VSS.n345 VSS.t133 5.8005
R3916 VSS.n345 VSS.t130 5.8005
R3917 VSS.n349 VSS.t35 5.8005
R3918 VSS.n349 VSS.t137 5.8005
R3919 VSS.n353 VSS.t28 5.8005
R3920 VSS.n353 VSS.t4 5.8005
R3921 VSS.n335 VSS.t29 5.8005
R3922 VSS.n335 VSS.t138 5.8005
R3923 VSS.n339 VSS.t132 5.8005
R3924 VSS.n339 VSS.t131 5.8005
R3925 VSS.n343 VSS.t58 5.8005
R3926 VSS.n343 VSS.t10 5.8005
R3927 VSS.n347 VSS.t134 5.8005
R3928 VSS.n347 VSS.t38 5.8005
R3929 VSS.n351 VSS.t42 5.8005
R3930 VSS.n351 VSS.t31 5.8005
R3931 VSS.n58 VSS.t56 5.8005
R3932 VSS.t86 VSS.n58 5.8005
R3933 VSS.n59 VSS.t86 5.8005
R3934 VSS.n59 VSS.t109 5.8005
R3935 VSS.n41 VSS.t2 5.8005
R3936 VSS.n41 VSS.t48 5.8005
R3937 VSS.n39 VSS.t46 5.8005
R3938 VSS.n39 VSS.t50 5.8005
R3939 VSS.n37 VSS.t34 5.8005
R3940 VSS.n37 VSS.t128 5.8005
R3941 VSS.n35 VSS.t8 5.8005
R3942 VSS.n35 VSS.t14 5.8005
R3943 VSS.n33 VSS.t55 5.8005
R3944 VSS.n33 VSS.t127 5.8005
R3945 VSS.n29 VSS.t118 5.8005
R3946 VSS.n29 VSS.t27 5.8005
R3947 VSS.n22 VSS.t120 5.8005
R3948 VSS.n22 VSS.t118 5.8005
R3949 VSS.n2302 VSS.t52 5.73102
R3950 VSS.n117 VSS.t36 5.73102
R3951 VSS.t5 VSS.t57 5.73102
R3952 VSS.t41 VSS.t59 5.73102
R3953 VSS.n285 VSS.n232 5.64756
R3954 VSS.n2513 VSS.n2503 5.64756
R3955 VSS.n66 VSS.n62 5.37662
R3956 VSS.n21 VSS.n9 5.37662
R3957 VSS.n1270 VSS.n1250 5.27109
R3958 VSS.n1215 VSS.n1203 5.27109
R3959 VSS.n1364 VSS.n1343 5.27109
R3960 VSS.n1858 VSS.n1857 5.27109
R3961 VSS.n1732 VSS.n1730 5.27109
R3962 VSS.n2101 VSS.n2100 5.27109
R3963 VSS.n2186 VSS.n2185 5.27109
R3964 VSS.n1178 VSS.n935 5.27109
R3965 VSS.t59 VSS.n1187 5.21007
R3966 VSS.n2095 VSS.t19 5.21007
R3967 VSS.n2296 VSS.n2295 4.68911
R3968 VSS.t41 VSS.n767 4.68911
R3969 VSS.n284 VSS.n234 4.51815
R3970 VSS.n397 VSS.n396 4.51815
R3971 VSS.n2517 VSS.n2502 4.51815
R3972 VSS.n2507 VSS.n76 4.51815
R3973 VSS.n1835 VSS.n1834 4.51815
R3974 VSS.n1885 VSS.n868 4.51815
R3975 VSS.n2179 VSS.n664 4.51815
R3976 VSS.n1953 VSS.n1952 4.51815
R3977 VSS.n1336 VSS.n885 4.5005
R3978 VSS.n1884 VSS.n1337 4.5005
R3979 VSS.n1888 VSS.n1887 4.5005
R3980 VSS.n1889 VSS.n866 4.5005
R3981 VSS.n1894 VSS.n1890 4.5005
R3982 VSS.n1899 VSS.n1898 4.5005
R3983 VSS.n1897 VSS.n1333 4.5005
R3984 VSS.n1896 VSS.n1895 4.5005
R3985 VSS.n1818 VSS.n1334 4.5005
R3986 VSS.n1392 VSS.n1391 4.5005
R3987 VSS.n1295 VSS.n1294 4.5005
R3988 VSS.n1296 VSS.n666 4.5005
R3989 VSS.n1911 VSS.n1297 4.5005
R3990 VSS.n1913 VSS.n1912 4.5005
R3991 VSS.n1915 VSS.n1914 4.5005
R3992 VSS.n1916 VSS.n1181 4.5005
R3993 VSS.n1948 VSS.n1180 4.5005
R3994 VSS.n1946 VSS.n1945 4.5005
R3995 VSS.n1947 VSS.n933 4.5005
R3996 VSS.n1950 VSS.n1949 4.5005
R3997 VSS.n2562 VSS.n73 4.26732
R3998 VSS.n2200 VSS.n527 4.22147
R3999 VSS.n1724 VSS.n1723 4.16815
R4000 VSS.n32 VSS.n3 3.81995
R4001 VSS.n326 VSS.n300 3.76521
R4002 VSS.n298 VSS.n296 3.76521
R4003 VSS.n303 VSS.n302 3.76521
R4004 VSS.n373 VSS.n371 3.76521
R4005 VSS.n386 VSS.n375 3.76521
R4006 VSS.n358 VSS.n357 3.76521
R4007 VSS.n69 VSS.n45 3.76521
R4008 VSS.n56 VSS.n50 3.76521
R4009 VSS.n28 VSS.n5 3.76521
R4010 VSS.n15 VSS.n14 3.76521
R4011 VSS.n1759 VSS.n1757 3.76521
R4012 VSS.n1274 VSS.n1273 3.76521
R4013 VSS.n1214 VSS.n1205 3.76521
R4014 VSS.n1365 VSS.n1341 3.76521
R4015 VSS.n1854 VSS.n1846 3.76521
R4016 VSS.n1819 VSS.n1816 3.76521
R4017 VSS.n2114 VSS.n867 3.76521
R4018 VSS.n2177 VSS.n665 3.76521
R4019 VSS.n1183 VSS.n930 3.76521
R4020 VSS.n2158 VSS.n698 3.76521
R4021 VSS.t5 VSS.n1904 3.6472
R4022 VSS.n2143 VSS.t23 3.6472
R4023 VSS.n2563 VSS.n2562 3.44797
R4024 VSS.n1257 VSS.n1255 3.09986
R4025 VSS.n1230 VSS.n1198 3.09986
R4026 VSS.n1351 VSS.n1350 3.09986
R4027 VSS.n1868 VSS.n1838 3.09986
R4028 VSS VSS.n2564 2.95131
R4029 VSS.n332 VSS.n331 2.89851
R4030 VSS.n376 VSS.n355 2.89851
R4031 VSS.n1336 VSS.n1335 2.78914
R4032 VSS.n1948 VSS.n527 2.78914
R4033 VSS.n51 VSS.n43 2.67025
R4034 VSS.n73 VSS.n72 2.67025
R4035 VSS.n32 VSS.n31 2.67025
R4036 VSS.n1822 VSS.n1821 2.63579
R4037 VSS.n2116 VSS.n865 2.63579
R4038 VSS.n2175 VSS.n667 2.63579
R4039 VSS.n1943 VSS.n1942 2.63579
R4040 VSS.n2071 VSS.n914 2.63579
R4041 VSS.n1427 VSS.t0 2.60528
R4042 VSS.n2103 VSS.t40 2.60528
R4043 VSS.n1335 VSS.n527 2.59582
R4044 VSS.t107 VSS.n1282 2.48621
R4045 VSS.n1282 VSS.t104 2.48621
R4046 VSS.t92 VSS.n1283 2.48621
R4047 VSS.n1283 VSS.t107 2.48621
R4048 VSS.t76 VSS.n1284 2.48621
R4049 VSS.n1284 VSS.t92 2.48621
R4050 VSS.t124 VSS.n1285 2.48621
R4051 VSS.n1285 VSS.t76 2.48621
R4052 VSS.n1231 VSS.t63 2.48621
R4053 VSS.t78 VSS.n1231 2.48621
R4054 VSS.n1232 VSS.t78 2.48621
R4055 VSS.t98 VSS.n1232 2.48621
R4056 VSS.n1233 VSS.t98 2.48621
R4057 VSS.t116 VSS.n1233 2.48621
R4058 VSS.n1234 VSS.t116 2.48621
R4059 VSS.t112 VSS.n1234 2.48621
R4060 VSS.n1286 VSS.t112 2.48621
R4061 VSS.n1286 VSS.t124 2.48621
R4062 VSS.t102 VSS.n1382 2.48621
R4063 VSS.n1382 VSS.t100 2.48621
R4064 VSS.t100 VSS.n1381 2.48621
R4065 VSS.n1381 VSS.t96 2.48621
R4066 VSS.t96 VSS.n1380 2.48621
R4067 VSS.n1380 VSS.t94 2.48621
R4068 VSS.t94 VSS.n1379 2.48621
R4069 VSS.n1379 VSS.t114 2.48621
R4070 VSS.t114 VSS.n1378 2.48621
R4071 VSS.n1378 VSS.t67 2.48621
R4072 VSS.t126 VSS.n1383 2.48621
R4073 VSS.n1383 VSS.t102 2.48621
R4074 VSS.t61 VSS.n1384 2.48621
R4075 VSS.n1384 VSS.t126 2.48621
R4076 VSS.t65 VSS.n1385 2.48621
R4077 VSS.n1385 VSS.t61 2.48621
R4078 VSS.n1872 VSS.t70 2.48621
R4079 VSS.n1872 VSS.t65 2.48621
R4080 VSS.n1391 VSS.n1390 2.30235
R4081 VSS.n1295 VSS.n659 2.30235
R4082 VSS.n307 VSS.n304 2.25932
R4083 VSS.n362 VSS.n359 2.25932
R4084 VSS.n68 VSS.n47 2.25932
R4085 VSS.n18 VSS.n10 2.25932
R4086 VSS.n1277 VSS.n1248 2.25932
R4087 VSS.n1211 VSS.n1210 2.25932
R4088 VSS.n1369 VSS.n1368 2.25932
R4089 VSS.n1853 VSS.n1848 2.25932
R4090 VSS.n315 VSS.n74 2.25177
R4091 VSS.n393 VSS.n392 2.25177
R4092 VSS.n2143 VSS.t21 2.08433
R4093 VSS.n2121 VSS.t17 2.08433
R4094 VSS.n1890 VSS.n1889 2.00152
R4095 VSS.n1898 VSS.n1334 2.00152
R4096 VSS.n1297 VSS.n1296 2.00152
R4097 VSS.n1946 VSS.n1181 2.00152
R4098 VSS.n1763 VSS.n1762 1.94348
R4099 VSS.n272 VSS.n271 1.88285
R4100 VSS.n281 VSS.n280 1.88285
R4101 VSS.n2528 VSS.n2499 1.88285
R4102 VSS.n2521 VSS.n2520 1.88285
R4103 VSS.n394 VSS.n393 1.82125
R4104 VSS.n2564 VSS.n2563 1.74238
R4105 VSS.n437 VSS.t83 1.56337
R4106 VSS.t72 VSS.n104 1.56337
R4107 VSS.t16 VSS.n673 1.56337
R4108 VSS.n2561 VSS.n2560 1.20384
R4109 VSS.n34 VSS.n32 1.1502
R4110 VSS.n36 VSS.n34 1.1502
R4111 VSS.n38 VSS.n36 1.1502
R4112 VSS.n40 VSS.n38 1.1502
R4113 VSS.n42 VSS.n40 1.1502
R4114 VSS.n43 VSS.n42 1.1502
R4115 VSS.n73 VSS.n43 1.1502
R4116 VSS.n1832 VSS.t6 1.04241
R4117 VSS.n2562 VSS.n2561 0.950967
R4118 VSS.n1281 VSS.n1280 0.779912
R4119 VSS.n1281 VSS.n1245 0.779912
R4120 VSS.n1245 VSS.n1244 0.779912
R4121 VSS.n1244 VSS.n1235 0.779912
R4122 VSS.n1291 VSS.n1196 0.779912
R4123 VSS.n1291 VSS.n1290 0.779912
R4124 VSS.n1290 VSS.n1289 0.779912
R4125 VSS.n1289 VSS.n1288 0.779912
R4126 VSS.n1288 VSS.n1287 0.779912
R4127 VSS.n1287 VSS.n1235 0.779912
R4128 VSS.n1877 VSS.n1375 0.779912
R4129 VSS.n1376 VSS.n1375 0.779912
R4130 VSS.n1377 VSS.n1376 0.779912
R4131 VSS.n1377 VSS.n1373 0.779912
R4132 VSS.n1373 VSS.n1372 0.779912
R4133 VSS.n1877 VSS.n1876 0.779912
R4134 VSS.n1876 VSS.n1875 0.779912
R4135 VSS.n1875 VSS.n1874 0.779912
R4136 VSS.n1873 VSS.n1386 0.779912
R4137 VSS.n1874 VSS.n1873 0.779912
R4138 VSS.n65 VSS.n64 0.753441
R4139 VSS.n20 VSS.n19 0.753441
R4140 VSS.n293 VSS.n292 0.753441
R4141 VSS.n2510 VSS.n2506 0.753441
R4142 VSS.n1761 VSS.n1760 0.753441
R4143 VSS.n1902 VSS.n1901 0.753441
R4144 VSS.n2145 VSS.n756 0.753441
R4145 VSS.n1909 VSS.n1908 0.753441
R4146 VSS.n1919 VSS.n1918 0.753441
R4147 VSS.n1239 VSS.n1238 0.701719
R4148 VSS.n1238 VSS.n1237 0.701719
R4149 VSS.n1237 VSS.n1236 0.701719
R4150 VSS.n1240 VSS.n1195 0.701719
R4151 VSS.n1241 VSS.n1240 0.701719
R4152 VSS.n1242 VSS.n1241 0.701719
R4153 VSS.n1880 VSS.n1879 0.701719
R4154 VSS.n1881 VSS.n1880 0.701719
R4155 VSS.n1882 VSS.n1881 0.701719
R4156 VSS.n1389 VSS.n1388 0.701719
R4157 VSS.n1388 VSS.n1387 0.701719
R4158 VSS.n1387 VSS.n1374 0.701719
R4159 VSS.n316 VSS.n315 0.647239
R4160 VSS.n392 VSS.n391 0.647239
R4161 VSS.n2561 VSS.n74 0.617976
R4162 VSS.n393 VSS.n355 0.574311
R4163 VSS.n355 VSS.n354 0.574311
R4164 VSS.n354 VSS.n352 0.574311
R4165 VSS.n352 VSS.n350 0.574311
R4166 VSS.n350 VSS.n348 0.574311
R4167 VSS.n348 VSS.n346 0.574311
R4168 VSS.n346 VSS.n344 0.574311
R4169 VSS.n344 VSS.n342 0.574311
R4170 VSS.n342 VSS.n340 0.574311
R4171 VSS.n340 VSS.n338 0.574311
R4172 VSS.n338 VSS.n336 0.574311
R4173 VSS.n336 VSS.n334 0.574311
R4174 VSS.n334 VSS.n332 0.574311
R4175 VSS.n332 VSS.n74 0.574311
R4176 VSS.n1335 VSS.n916 0.538331
R4177 VSS.n2347 VSS.t7 0.521457
R4178 VSS.n2408 VSS.t11 0.521457
R4179 VSS.n315 VSS.n314 0.418978
R4180 VSS.n392 VSS.n369 0.418978
R4181 VSS.n320 VSS.n319 0.320353
R4182 VSS.n322 VSS.n320 0.320353
R4183 VSS.n322 VSS.n321 0.320353
R4184 VSS.n306 VSS.n305 0.320353
R4185 VSS.n382 VSS.n381 0.320353
R4186 VSS.n380 VSS.n377 0.320353
R4187 VSS.n381 VSS.n380 0.320353
R4188 VSS.n361 VSS.n360 0.320353
R4189 VSS.n52 VSS.n48 0.320353
R4190 VSS.n60 VSS.n48 0.320353
R4191 VSS.n61 VSS.n60 0.320353
R4192 VSS.n66 VSS.n61 0.320353
R4193 VSS.n9 VSS.n7 0.320353
R4194 VSS.n23 VSS.n7 0.320353
R4195 VSS.n24 VSS.n23 0.320353
R4196 VSS.n25 VSS.n24 0.320353
R4197 VSS.n2563 VSS.n2 0.303278
R4198 VSS.n2564 VSS.n1 0.303278
R4199 VSS.n1281 VSS.n932 0.272321
R4200 VSS.n1292 VSS.n1291 0.272321
R4201 VSS.n1287 VSS.n1243 0.272321
R4202 VSS.n1883 VSS.n1373 0.272321
R4203 VSS.n1878 VSS.n1877 0.272321
R4204 VSS.n1873 VSS.n1837 0.272321
R4205 VSS.n1243 VSS.n1239 0.261436
R4206 VSS.n1236 VSS.n932 0.261436
R4207 VSS.n1292 VSS.n1195 0.261436
R4208 VSS.n1243 VSS.n1242 0.261436
R4209 VSS.n1879 VSS.n1878 0.261436
R4210 VSS.n1883 VSS.n1882 0.261436
R4211 VSS.n1837 VSS.n1389 0.261436
R4212 VSS.n1878 VSS.n1374 0.261436
R4213 VSS VSS.n0 0.245958
R4214 VSS.n2523 VSS.n2522 0.243804
R4215 VSS.n2512 VSS.n2501 0.243804
R4216 VSS.n282 VSS.n235 0.243804
R4217 VSS.n283 VSS.n231 0.243804
R4218 VSS.n2200 VSS.n2199 0.21925
R4219 VSS.n2511 VSS.n75 0.204927
R4220 VSS.n395 VSS.n294 0.204927
R4221 VSS.n835 VSS.n832 0.204369
R4222 VSS.n847 VSS.n846 0.204369
R4223 VSS.n331 VSS.n295 0.196152
R4224 VSS.n318 VSS.n295 0.196152
R4225 VSS.n319 VSS.n318 0.196152
R4226 VSS.n309 VSS.n306 0.196152
R4227 VSS.n309 VSS.n308 0.196152
R4228 VSS.n308 VSS.n301 0.196152
R4229 VSS.n314 VSS.n301 0.196152
R4230 VSS.n325 VSS.n316 0.196152
R4231 VSS.n325 VSS.n324 0.196152
R4232 VSS.n324 VSS.n322 0.196152
R4233 VSS.n385 VSS.n376 0.196152
R4234 VSS.n385 VSS.n384 0.196152
R4235 VSS.n384 VSS.n382 0.196152
R4236 VSS.n364 VSS.n361 0.196152
R4237 VSS.n364 VSS.n363 0.196152
R4238 VSS.n363 VSS.n356 0.196152
R4239 VSS.n369 VSS.n356 0.196152
R4240 VSS.n391 VSS.n370 0.196152
R4241 VSS.n379 VSS.n370 0.196152
R4242 VSS.n380 VSS.n379 0.196152
R4243 VSS.n55 VSS.n51 0.196152
R4244 VSS.n55 VSS.n54 0.196152
R4245 VSS.n54 VSS.n52 0.196152
R4246 VSS.n72 VSS.n44 0.196152
R4247 VSS.n67 VSS.n44 0.196152
R4248 VSS.n67 VSS.n66 0.196152
R4249 VSS.n13 VSS.n3 0.196152
R4250 VSS.n13 VSS.n12 0.196152
R4251 VSS.n12 VSS.n9 0.196152
R4252 VSS.n31 VSS.n4 0.196152
R4253 VSS.n26 VSS.n4 0.196152
R4254 VSS.n26 VSS.n25 0.196152
R4255 VSS.n1280 VSS.n1279 0.196152
R4256 VSS.n1279 VSS.n1247 0.196152
R4257 VSS.n1272 VSS.n1247 0.196152
R4258 VSS.n1272 VSS.n1271 0.196152
R4259 VSS.n1271 VSS.n1251 0.196152
R4260 VSS.n1264 VSS.n1251 0.196152
R4261 VSS.n1264 VSS.n1263 0.196152
R4262 VSS.n1263 VSS.n1255 0.196152
R4263 VSS.n1206 VSS.n1196 0.196152
R4264 VSS.n1212 VSS.n1206 0.196152
R4265 VSS.n1213 VSS.n1212 0.196152
R4266 VSS.n1213 VSS.n1202 0.196152
R4267 VSS.n1220 VSS.n1202 0.196152
R4268 VSS.n1222 VSS.n1220 0.196152
R4269 VSS.n1222 VSS.n1221 0.196152
R4270 VSS.n1221 VSS.n1198 0.196152
R4271 VSS.n1351 VSS.n1346 0.196152
R4272 VSS.n1358 VSS.n1346 0.196152
R4273 VSS.n1359 VSS.n1358 0.196152
R4274 VSS.n1359 VSS.n1342 0.196152
R4275 VSS.n1366 VSS.n1342 0.196152
R4276 VSS.n1367 VSS.n1366 0.196152
R4277 VSS.n1367 VSS.n1338 0.196152
R4278 VSS.n1372 VSS.n1338 0.196152
R4279 VSS.n1868 VSS.n1867 0.196152
R4280 VSS.n1867 VSS.n1841 0.196152
R4281 VSS.n1860 VSS.n1841 0.196152
R4282 VSS.n1860 VSS.n1859 0.196152
R4283 VSS.n1859 VSS.n1845 0.196152
R4284 VSS.n1852 VSS.n1845 0.196152
R4285 VSS.n1852 VSS.n1851 0.196152
R4286 VSS.n1851 VSS.n1386 0.196152
R4287 VSS.n2522 VSS.n2501 0.190232
R4288 VSS.n2512 VSS.n2511 0.190232
R4289 VSS.n283 VSS.n282 0.190232
R4290 VSS.n294 VSS.n231 0.190232
R4291 VSS.n1950 VSS.n1180 0.146333
R4292 VSS.n1945 VSS.n933 0.146333
R4293 VSS.n1916 VSS.n1915 0.146333
R4294 VSS.n1912 VSS.n1911 0.146333
R4295 VSS.n1899 VSS.n1333 0.146333
R4296 VSS.n1895 VSS.n1894 0.146333
R4297 VSS.n1887 VSS.n866 0.146333
R4298 VSS.n1884 VSS.n885 0.146333
R4299 VSS.n1818 VSS.n1392 0.146333
R4300 VSS.n1294 VSS.n666 0.146333
R4301 VSS.n1731 VSS.n1390 0.144812
R4302 VSS.n2187 VSS.n659 0.144812
R4303 VSS.n1836 VSS.n1390 0.119763
R4304 VSS.n1293 VSS.n659 0.119763
R4305 VSS.n846 VSS.n832 0.119548
R4306 VSS.n1951 VSS.n932 0.114136
R4307 VSS.n1293 VSS.n1292 0.114136
R4308 VSS.n1243 VSS.n1194 0.114136
R4309 VSS.n1886 VSS.n1883 0.114136
R4310 VSS.n1878 VSS.n755 0.114136
R4311 VSS.n1837 VSS.n1836 0.114136
R4312 VSS.n1756 VSS.n1755 0.113595
R4313 VSS.n2560 VSS.n75 0.104667
R4314 VSS.n395 VSS.n394 0.104667
R4315 VSS.n1889 VSS.n1888 0.0788898
R4316 VSS.n1337 VSS.n1336 0.0788898
R4317 VSS.n1898 VSS.n1897 0.0788898
R4318 VSS.n1896 VSS.n1890 0.0788898
R4319 VSS.n1391 VSS.n1334 0.0788898
R4320 VSS.n1296 VSS.n1295 0.0788898
R4321 VSS.n1913 VSS.n1297 0.0788898
R4322 VSS.n1914 VSS.n1181 0.0788898
R4323 VSS.n1947 VSS.n1946 0.0788898
R4324 VSS.n1949 VSS.n1948 0.0788898
R4325 VSS.n1180 VSS.n1179 0.0719286
R4326 VSS.n1945 VSS.n1944 0.0719286
R4327 VSS.n1917 VSS.n1916 0.0719286
R4328 VSS.n1911 VSS.n1910 0.0719286
R4329 VSS.n1900 VSS.n1899 0.0719286
R4330 VSS.n1894 VSS.n1893 0.0719286
R4331 VSS.n2115 VSS.n866 0.0719286
R4332 VSS.n2099 VSS.n885 0.0719286
R4333 VSS.n1820 VSS.n1818 0.0719286
R4334 VSS.n2176 VSS.n666 0.0719286
R4335 VSS.n1888 VSS.n1337 0.0682966
R4336 VSS.n1897 VSS.n1896 0.0682966
R4337 VSS.n1914 VSS.n1913 0.0682966
R4338 VSS.n1949 VSS.n1947 0.0682966
R4339 VSS.n847 VSS.n1 0.0615119
R4340 VSS.n1756 VSS.n2 0.0600238
R4341 VSS.n1762 VSS.n2 0.0600238
R4342 VSS.n1951 VSS.n933 0.048119
R4343 VSS.n1951 VSS.n1950 0.048119
R4344 VSS.n1912 VSS.n1194 0.048119
R4345 VSS.n1915 VSS.n1194 0.048119
R4346 VSS.n1333 VSS.n755 0.048119
R4347 VSS.n1895 VSS.n755 0.048119
R4348 VSS.n1887 VSS.n1886 0.048119
R4349 VSS.n1886 VSS.n1884 0.048119
R4350 VSS.n1836 VSS.n1392 0.048119
R4351 VSS.n1294 VSS.n1293 0.048119
R4352 VSS.n2066 VSS.n2065 0.0344109
R4353 VSS.n922 VSS.n917 0.0344109
R4354 VSS.n2066 VSS.n916 0.020302
R4355 VSS.n2065 VSS.n917 0.020302
R4356 VSS.n922 VSS.n0 0.020302
R4357 a_2479_7336.n0 a_2479_7336.t31 260.486
R4358 a_2479_7336.n68 a_2479_7336.t19 260.486
R4359 a_2479_7336.n79 a_2479_7336.t34 260.111
R4360 a_2479_7336.n80 a_2479_7336.t21 260.111
R4361 a_2479_7336.n81 a_2479_7336.t29 260.111
R4362 a_2479_7336.n82 a_2479_7336.t18 260.111
R4363 a_2479_7336.n83 a_2479_7336.t33 260.111
R4364 a_2479_7336.n84 a_2479_7336.t27 260.111
R4365 a_2479_7336.n1 a_2479_7336.t24 260.111
R4366 a_2479_7336.n0 a_2479_7336.t22 260.111
R4367 a_2479_7336.n68 a_2479_7336.t28 260.111
R4368 a_2479_7336.n69 a_2479_7336.t35 260.111
R4369 a_2479_7336.n71 a_2479_7336.t32 260.111
R4370 a_2479_7336.n72 a_2479_7336.t26 260.111
R4371 a_2479_7336.n73 a_2479_7336.t23 260.111
R4372 a_2479_7336.n74 a_2479_7336.t20 260.111
R4373 a_2479_7336.n75 a_2479_7336.t30 260.111
R4374 a_2479_7336.n76 a_2479_7336.t25 260.111
R4375 a_2479_7336.n86 a_2479_7336.n85 203.843
R4376 a_2479_7336.n70 a_2479_7336.n67 203.843
R4377 a_2479_7336.n59 a_2479_7336.n41 185
R4378 a_2479_7336.n59 a_2479_7336.n40 185
R4379 a_2479_7336.n59 a_2479_7336.n39 185
R4380 a_2479_7336.n59 a_2479_7336.n38 185
R4381 a_2479_7336.n59 a_2479_7336.n37 185
R4382 a_2479_7336.n59 a_2479_7336.n36 185
R4383 a_2479_7336.n59 a_2479_7336.n35 185
R4384 a_2479_7336.n28 a_2479_7336.n10 185
R4385 a_2479_7336.n28 a_2479_7336.n9 185
R4386 a_2479_7336.n28 a_2479_7336.n8 185
R4387 a_2479_7336.n28 a_2479_7336.n7 185
R4388 a_2479_7336.n28 a_2479_7336.n6 185
R4389 a_2479_7336.n28 a_2479_7336.n5 185
R4390 a_2479_7336.n28 a_2479_7336.n4 185
R4391 a_2479_7336.n43 a_2479_7336.t11 130.75
R4392 a_2479_7336.n12 a_2479_7336.t14 130.75
R4393 a_2479_7336.n43 a_2479_7336.t13 91.3557
R4394 a_2479_7336.n12 a_2479_7336.t15 91.3557
R4395 a_2479_7336.n60 a_2479_7336.n59 86.5152
R4396 a_2479_7336.n29 a_2479_7336.n28 86.5152
R4397 a_2479_7336.n58 a_2479_7336.n42 30.3012
R4398 a_2479_7336.n27 a_2479_7336.n11 30.3012
R4399 a_2479_7336.n67 a_2479_7336.t10 28.5655
R4400 a_2479_7336.n67 a_2479_7336.t8 28.5655
R4401 a_2479_7336.t0 a_2479_7336.n86 28.5655
R4402 a_2479_7336.n86 a_2479_7336.t2 28.5655
R4403 a_2479_7336.n35 a_2479_7336.n34 24.8476
R4404 a_2479_7336.n4 a_2479_7336.n3 24.8476
R4405 a_2479_7336.n44 a_2479_7336.n36 23.3417
R4406 a_2479_7336.n13 a_2479_7336.n5 23.3417
R4407 a_2479_7336.n61 a_2479_7336.n60 22.0256
R4408 a_2479_7336.n30 a_2479_7336.n29 22.0256
R4409 a_2479_7336.n46 a_2479_7336.n37 21.8358
R4410 a_2479_7336.n15 a_2479_7336.n6 21.8358
R4411 a_2479_7336.n48 a_2479_7336.n38 20.3299
R4412 a_2479_7336.n17 a_2479_7336.n7 20.3299
R4413 a_2479_7336.n50 a_2479_7336.n39 18.824
R4414 a_2479_7336.n19 a_2479_7336.n8 18.824
R4415 a_2479_7336.n52 a_2479_7336.n40 17.3181
R4416 a_2479_7336.n21 a_2479_7336.n9 17.3181
R4417 a_2479_7336.n59 a_2479_7336.n58 16.3559
R4418 a_2479_7336.n28 a_2479_7336.n27 16.3559
R4419 a_2479_7336.n54 a_2479_7336.n41 15.8123
R4420 a_2479_7336.n23 a_2479_7336.n10 15.8123
R4421 a_2479_7336.n64 a_2479_7336.n63 14.6052
R4422 a_2479_7336.n66 a_2479_7336.n65 14.6052
R4423 a_2479_7336.n32 a_2479_7336.n31 14.377
R4424 a_2479_7336.n60 a_2479_7336.n34 12.7256
R4425 a_2479_7336.n29 a_2479_7336.n3 12.7256
R4426 a_2479_7336.n77 a_2479_7336.t9 12.5928
R4427 a_2479_7336.n64 a_2479_7336.n62 11.5586
R4428 a_2479_7336.n42 a_2479_7336.n41 11.2946
R4429 a_2479_7336.n11 a_2479_7336.n10 11.2946
R4430 a_2479_7336.n54 a_2479_7336.n40 9.78874
R4431 a_2479_7336.n23 a_2479_7336.n9 9.78874
R4432 a_2479_7336.n34 a_2479_7336.n33 9.3005
R4433 a_2479_7336.n45 a_2479_7336.n44 9.3005
R4434 a_2479_7336.n47 a_2479_7336.n46 9.3005
R4435 a_2479_7336.n49 a_2479_7336.n48 9.3005
R4436 a_2479_7336.n51 a_2479_7336.n50 9.3005
R4437 a_2479_7336.n53 a_2479_7336.n52 9.3005
R4438 a_2479_7336.n55 a_2479_7336.n54 9.3005
R4439 a_2479_7336.n56 a_2479_7336.n42 9.3005
R4440 a_2479_7336.n3 a_2479_7336.n2 9.3005
R4441 a_2479_7336.n14 a_2479_7336.n13 9.3005
R4442 a_2479_7336.n16 a_2479_7336.n15 9.3005
R4443 a_2479_7336.n18 a_2479_7336.n17 9.3005
R4444 a_2479_7336.n20 a_2479_7336.n19 9.3005
R4445 a_2479_7336.n22 a_2479_7336.n21 9.3005
R4446 a_2479_7336.n24 a_2479_7336.n23 9.3005
R4447 a_2479_7336.n25 a_2479_7336.n11 9.3005
R4448 a_2479_7336.n52 a_2479_7336.n39 8.28285
R4449 a_2479_7336.n21 a_2479_7336.n8 8.28285
R4450 a_2479_7336.n78 a_2479_7336.n66 8.22405
R4451 a_2479_7336.n50 a_2479_7336.n38 6.77697
R4452 a_2479_7336.n19 a_2479_7336.n7 6.77697
R4453 a_2479_7336.n32 a_2479_7336.n30 6.19091
R4454 a_2479_7336.n48 a_2479_7336.n37 5.27109
R4455 a_2479_7336.n17 a_2479_7336.n6 5.27109
R4456 a_2479_7336.n78 a_2479_7336.n77 4.66982
R4457 a_2479_7336.n46 a_2479_7336.n36 3.76521
R4458 a_2479_7336.n15 a_2479_7336.n5 3.76521
R4459 a_2479_7336.n62 a_2479_7336.n61 3.31388
R4460 a_2479_7336.n66 a_2479_7336.n64 2.87753
R4461 a_2479_7336.n63 a_2479_7336.t16 2.48621
R4462 a_2479_7336.n63 a_2479_7336.t17 2.48621
R4463 a_2479_7336.n65 a_2479_7336.t4 2.48621
R4464 a_2479_7336.n65 a_2479_7336.t3 2.48621
R4465 a_2479_7336.n59 a_2479_7336.t5 2.48621
R4466 a_2479_7336.n59 a_2479_7336.t12 2.48621
R4467 a_2479_7336.n28 a_2479_7336.t15 2.48621
R4468 a_2479_7336.n28 a_2479_7336.t6 2.48621
R4469 a_2479_7336.n31 a_2479_7336.t1 2.48621
R4470 a_2479_7336.n31 a_2479_7336.t7 2.48621
R4471 a_2479_7336.n58 a_2479_7336.n57 2.36936
R4472 a_2479_7336.n27 a_2479_7336.n26 2.36936
R4473 a_2479_7336.n62 a_2479_7336.n32 2.30287
R4474 a_2479_7336.n44 a_2479_7336.n35 2.25932
R4475 a_2479_7336.n13 a_2479_7336.n4 2.25932
R4476 a_2479_7336.n77 a_2479_7336.n76 1.41083
R4477 a_2479_7336.n79 a_2479_7336.n78 1.3088
R4478 a_2479_7336.n76 a_2479_7336.n75 0.3755
R4479 a_2479_7336.n75 a_2479_7336.n74 0.3755
R4480 a_2479_7336.n74 a_2479_7336.n73 0.3755
R4481 a_2479_7336.n73 a_2479_7336.n72 0.3755
R4482 a_2479_7336.n72 a_2479_7336.n71 0.3755
R4483 a_2479_7336.n69 a_2479_7336.n68 0.3755
R4484 a_2479_7336.n1 a_2479_7336.n0 0.3755
R4485 a_2479_7336.n84 a_2479_7336.n83 0.3755
R4486 a_2479_7336.n83 a_2479_7336.n82 0.3755
R4487 a_2479_7336.n82 a_2479_7336.n81 0.3755
R4488 a_2479_7336.n81 a_2479_7336.n80 0.3755
R4489 a_2479_7336.n80 a_2479_7336.n79 0.3755
R4490 a_2479_7336.n57 a_2479_7336.n43 0.320353
R4491 a_2479_7336.n26 a_2479_7336.n12 0.320353
R4492 a_2479_7336.n57 a_2479_7336.n56 0.196152
R4493 a_2479_7336.n56 a_2479_7336.n55 0.196152
R4494 a_2479_7336.n55 a_2479_7336.n53 0.196152
R4495 a_2479_7336.n53 a_2479_7336.n51 0.196152
R4496 a_2479_7336.n51 a_2479_7336.n49 0.196152
R4497 a_2479_7336.n49 a_2479_7336.n47 0.196152
R4498 a_2479_7336.n47 a_2479_7336.n45 0.196152
R4499 a_2479_7336.n45 a_2479_7336.n33 0.196152
R4500 a_2479_7336.n61 a_2479_7336.n33 0.196152
R4501 a_2479_7336.n26 a_2479_7336.n25 0.196152
R4502 a_2479_7336.n25 a_2479_7336.n24 0.196152
R4503 a_2479_7336.n24 a_2479_7336.n22 0.196152
R4504 a_2479_7336.n22 a_2479_7336.n20 0.196152
R4505 a_2479_7336.n20 a_2479_7336.n18 0.196152
R4506 a_2479_7336.n18 a_2479_7336.n16 0.196152
R4507 a_2479_7336.n16 a_2479_7336.n14 0.196152
R4508 a_2479_7336.n14 a_2479_7336.n2 0.196152
R4509 a_2479_7336.n30 a_2479_7336.n2 0.196152
R4510 a_2479_7336.n71 a_2479_7336.n70 0.188
R4511 a_2479_7336.n70 a_2479_7336.n69 0.188
R4512 a_2479_7336.n85 a_2479_7336.n1 0.188
R4513 a_2479_7336.n85 a_2479_7336.n84 0.188
R4514 VOUT.n13 VOUT.t8 260.298
R4515 VOUT.t4 VOUT.n13 260.298
R4516 VOUT.t8 VOUT.n8 260.298
R4517 VOUT.n56 VOUT.t6 260.298
R4518 VOUT.t2 VOUT.n56 260.298
R4519 VOUT.n57 VOUT.t2 260.298
R4520 VOUT.n14 VOUT.t4 260.111
R4521 VOUT.t6 VOUT.n54 260.111
R4522 VOUT.n12 VOUT.t10 232.03
R4523 VOUT.t3 VOUT.n55 232.03
R4524 VOUT.n2 VOUT.n0 206.708
R4525 VOUT.n6 VOUT.n5 206.094
R4526 VOUT.n4 VOUT.n3 206.094
R4527 VOUT.n2 VOUT.n1 206.094
R4528 VOUT.n70 VOUT.n69 206.094
R4529 VOUT.n68 VOUT.n67 206.094
R4530 VOUT.n66 VOUT.n65 206.094
R4531 VOUT.n64 VOUT.n63 206.094
R4532 VOUT.n11 VOUT.n10 203.03
R4533 VOUT.n9 VOUT.n7 203.03
R4534 VOUT.n61 VOUT.n60 203.03
R4535 VOUT.n59 VOUT.n58 203.03
R4536 VOUT.n43 VOUT.n42 185
R4537 VOUT.n43 VOUT.n25 185
R4538 VOUT.n43 VOUT.n24 185
R4539 VOUT.n43 VOUT.n23 185
R4540 VOUT.n43 VOUT.n22 185
R4541 VOUT.n43 VOUT.n21 185
R4542 VOUT.n43 VOUT.n20 185
R4543 VOUT.n26 VOUT.t11 130.75
R4544 VOUT.n26 VOUT.t13 91.3557
R4545 VOUT.n44 VOUT.n43 86.5152
R4546 VOUT.n28 VOUT.n19 30.3012
R4547 VOUT.n10 VOUT.t5 28.5655
R4548 VOUT.n10 VOUT.t9 28.5655
R4549 VOUT.n9 VOUT.t18 28.5655
R4550 VOUT.t5 VOUT.n9 28.5655
R4551 VOUT.n5 VOUT.t20 28.5655
R4552 VOUT.n5 VOUT.t17 28.5655
R4553 VOUT.n3 VOUT.t19 28.5655
R4554 VOUT.n3 VOUT.t14 28.5655
R4555 VOUT.n1 VOUT.t21 28.5655
R4556 VOUT.n1 VOUT.t16 28.5655
R4557 VOUT.n0 VOUT.t26 28.5655
R4558 VOUT.n0 VOUT.t28 28.5655
R4559 VOUT.n60 VOUT.t7 28.5655
R4560 VOUT.n60 VOUT.t22 28.5655
R4561 VOUT.n59 VOUT.t3 28.5655
R4562 VOUT.t7 VOUT.n59 28.5655
R4563 VOUT.n69 VOUT.t24 28.5655
R4564 VOUT.n69 VOUT.t27 28.5655
R4565 VOUT.n67 VOUT.t25 28.5655
R4566 VOUT.n67 VOUT.t15 28.5655
R4567 VOUT.n65 VOUT.t29 28.5655
R4568 VOUT.n65 VOUT.t31 28.5655
R4569 VOUT.n63 VOUT.t23 28.5655
R4570 VOUT.n63 VOUT.t30 28.5655
R4571 VOUT.n42 VOUT.n18 24.8476
R4572 VOUT.n41 VOUT.n25 23.3417
R4573 VOUT.n45 VOUT.n44 22.0256
R4574 VOUT.n38 VOUT.n24 21.8358
R4575 VOUT.n36 VOUT.n23 20.3299
R4576 VOUT.n46 VOUT.n45 19.0885
R4577 VOUT.n34 VOUT.n22 18.824
R4578 VOUT.n32 VOUT.n21 17.3181
R4579 VOUT.n43 VOUT.n19 16.3559
R4580 VOUT.n30 VOUT.n20 15.8123
R4581 VOUT.n44 VOUT.n18 12.7256
R4582 VOUT.n28 VOUT.n20 11.2946
R4583 VOUT.n30 VOUT.n21 9.78874
R4584 VOUT.n18 VOUT.n17 9.3005
R4585 VOUT.n41 VOUT.n40 9.3005
R4586 VOUT.n39 VOUT.n38 9.3005
R4587 VOUT.n37 VOUT.n36 9.3005
R4588 VOUT.n35 VOUT.n34 9.3005
R4589 VOUT.n33 VOUT.n32 9.3005
R4590 VOUT.n31 VOUT.n30 9.3005
R4591 VOUT.n29 VOUT.n28 9.3005
R4592 VOUT.n32 VOUT.n22 8.28285
R4593 VOUT.n34 VOUT.n23 6.77697
R4594 VOUT.n36 VOUT.n24 5.27109
R4595 VOUT.n38 VOUT.n25 3.76521
R4596 VOUT.n48 VOUT.n47 3.4105
R4597 VOUT.n72 VOUT.n46 3.29996
R4598 VOUT.n64 VOUT.n62 3.23261
R4599 VOUT.n16 VOUT.n15 2.55612
R4600 VOUT.n43 VOUT.t0 2.48621
R4601 VOUT.n43 VOUT.t12 2.48621
R4602 VOUT VOUT.n16 2.47337
R4603 VOUT.n27 VOUT.n19 2.36936
R4604 VOUT.n42 VOUT.n41 2.25932
R4605 VOUT.n71 VOUT.n70 2.12962
R4606 VOUT.n53 VOUT.n52 1.70927
R4607 VOUT.n51 VOUT.n50 1.7055
R4608 VOUT.n50 VOUT.n49 1.7055
R4609 VOUT.n52 VOUT.n51 1.14963
R4610 VOUT.n72 VOUT.n71 1.09816
R4611 VOUT.n4 VOUT.n2 0.61449
R4612 VOUT.n6 VOUT.n4 0.61449
R4613 VOUT.n16 VOUT.n6 0.61449
R4614 VOUT.n66 VOUT.n64 0.61449
R4615 VOUT.n68 VOUT.n66 0.61449
R4616 VOUT.n70 VOUT.n68 0.61449
R4617 VOUT.n51 VOUT.t1 0.563396
R4618 VOUT VOUT.n72 0.521984
R4619 VOUT.n62 VOUT.n61 0.446229
R4620 VOUT.n61 VOUT.n55 0.43664
R4621 VOUT.n12 VOUT.n7 0.436638
R4622 VOUT.n15 VOUT.n7 0.38373
R4623 VOUT.n11 VOUT.n8 0.38373
R4624 VOUT.n58 VOUT.n57 0.383729
R4625 VOUT.n27 VOUT.n26 0.320353
R4626 VOUT.n13 VOUT.n12 0.285826
R4627 VOUT.n56 VOUT.n55 0.285826
R4628 VOUT.n49 VOUT.n46 0.2193
R4629 VOUT.n45 VOUT.n17 0.196152
R4630 VOUT.n40 VOUT.n17 0.196152
R4631 VOUT.n40 VOUT.n39 0.196152
R4632 VOUT.n39 VOUT.n37 0.196152
R4633 VOUT.n37 VOUT.n35 0.196152
R4634 VOUT.n35 VOUT.n33 0.196152
R4635 VOUT.n33 VOUT.n31 0.196152
R4636 VOUT.n31 VOUT.n29 0.196152
R4637 VOUT.n29 VOUT.n27 0.196152
R4638 VOUT.n15 VOUT.n14 0.188
R4639 VOUT.n14 VOUT.n8 0.188
R4640 VOUT.n57 VOUT.n54 0.188
R4641 VOUT.n62 VOUT.n54 0.1255
R4642 VOUT.n58 VOUT.n55 0.0984044
R4643 VOUT.n12 VOUT.n11 0.0984028
R4644 VOUT.n71 VOUT.n53 0.0647077
R4645 VOUT.n50 VOUT.n48 0.0102917
R4646 VOUT.n52 VOUT.n48 0.00750288
R4647 VOUT.n53 VOUT.n47 0.00118306
R4648 VOUT.n49 VOUT.n47 0.00118306
R4649 VDD.n312 VDD.n67 723.529
R4650 VDD.n72 VDD.n64 723.529
R4651 VDD.n139 VDD.n111 723.529
R4652 VDD.n187 VDD.n113 723.529
R4653 VDD.n266 VDD.n265 515.294
R4654 VDD.n301 VDD.n52 275.295
R4655 VDD.n152 VDD.n132 275.295
R4656 VDD.n34 VDD.t54 260.486
R4657 VDD.n20 VDD.t29 260.486
R4658 VDD.n346 VDD.t18 260.486
R4659 VDD.n331 VDD.t38 260.486
R4660 VDD.t11 VDD.n38 260.298
R4661 VDD.n36 VDD.t32 260.298
R4662 VDD.n39 VDD.t11 260.298
R4663 VDD.t51 VDD.n19 260.298
R4664 VDD.n17 VDD.t40 260.298
R4665 VDD.n13 VDD.t40 260.298
R4666 VDD.t24 VDD.n343 260.298
R4667 VDD.t42 VDD.n345 260.298
R4668 VDD.n350 VDD.t24 260.298
R4669 VDD.n328 VDD.t49 260.298
R4670 VDD.t49 VDD.n325 260.298
R4671 VDD.n332 VDD.t56 260.298
R4672 VDD.n1 VDD.t21 260.199
R4673 VDD.n368 VDD.t44 260.199
R4674 VDD.t35 VDD.n32 260.111
R4675 VDD.n37 VDD.t35 260.111
R4676 VDD.t32 VDD.n34 260.111
R4677 VDD.n20 VDD.t51 260.111
R4678 VDD.t15 VDD.n12 260.111
R4679 VDD.n18 VDD.t15 260.111
R4680 VDD.n349 VDD.t47 260.111
R4681 VDD.t47 VDD.n348 260.111
R4682 VDD.n346 VDD.t42 260.111
R4683 VDD.t56 VDD.n331 260.111
R4684 VDD.n330 VDD.t27 260.111
R4685 VDD.t27 VDD.n329 260.111
R4686 VDD.n66 VDD.n65 240
R4687 VDD.n299 VDD.n65 240
R4688 VDD.n305 VDD.n304 240
R4689 VDD.n316 VDD.n51 240
R4690 VDD.n262 VDD.n261 240
R4691 VDD.n270 VDD.n269 240
R4692 VDD.n274 VDD.n273 240
R4693 VDD.n278 VDD.n277 240
R4694 VDD.n282 VDD.n281 240
R4695 VDD.n286 VDD.n285 240
R4696 VDD.n288 VDD.n64 240
R4697 VDD.n193 VDD.n111 240
R4698 VDD.n193 VDD.n109 240
R4699 VDD.n197 VDD.n109 240
R4700 VDD.n197 VDD.n104 240
R4701 VDD.n206 VDD.n104 240
R4702 VDD.n206 VDD.n102 240
R4703 VDD.n210 VDD.n102 240
R4704 VDD.n210 VDD.n97 240
R4705 VDD.n219 VDD.n97 240
R4706 VDD.n219 VDD.n95 240
R4707 VDD.n223 VDD.n95 240
R4708 VDD.n223 VDD.n90 240
R4709 VDD.n231 VDD.n90 240
R4710 VDD.n231 VDD.n88 240
R4711 VDD.n235 VDD.n88 240
R4712 VDD.n235 VDD.n82 240
R4713 VDD.n243 VDD.n82 240
R4714 VDD.n243 VDD.n80 240
R4715 VDD.n247 VDD.n80 240
R4716 VDD.n247 VDD.n74 240
R4717 VDD.n255 VDD.n74 240
R4718 VDD.n255 VDD.n71 240
R4719 VDD.n293 VDD.n71 240
R4720 VDD.n293 VDD.n72 240
R4721 VDD.n185 VDD.n184 240
R4722 VDD.n182 VDD.n118 240
R4723 VDD.n178 VDD.n177 240
R4724 VDD.n175 VDD.n121 240
R4725 VDD.n169 VDD.n168 240
R4726 VDD.n166 VDD.n126 240
R4727 VDD.n162 VDD.n161 240
R4728 VDD.n159 VDD.n129 240
R4729 VDD.n155 VDD.n154 240
R4730 VDD.n146 VDD.n145 240
R4731 VDD.n143 VDD.n137 240
R4732 VDD.n191 VDD.n113 240
R4733 VDD.n191 VDD.n108 240
R4734 VDD.n200 VDD.n108 240
R4735 VDD.n200 VDD.n106 240
R4736 VDD.n204 VDD.n106 240
R4737 VDD.n204 VDD.n101 240
R4738 VDD.n213 VDD.n101 240
R4739 VDD.n213 VDD.n99 240
R4740 VDD.n217 VDD.n99 240
R4741 VDD.n217 VDD.n94 240
R4742 VDD.n225 VDD.n94 240
R4743 VDD.n225 VDD.n92 240
R4744 VDD.n229 VDD.n92 240
R4745 VDD.n229 VDD.n86 240
R4746 VDD.n237 VDD.n86 240
R4747 VDD.n237 VDD.n84 240
R4748 VDD.n241 VDD.n84 240
R4749 VDD.n241 VDD.n78 240
R4750 VDD.n249 VDD.n78 240
R4751 VDD.n249 VDD.n76 240
R4752 VDD.n253 VDD.n76 240
R4753 VDD.n253 VDD.n69 240
R4754 VDD.n295 VDD.n69 240
R4755 VDD.n295 VDD.n67 240
R4756 VDD.n31 VDD.t14 232.03
R4757 VDD.n16 VDD.t41 232.03
R4758 VDD.n351 VDD.t26 232.03
R4759 VDD.t50 VDD.n324 232.03
R4760 VDD.n367 VDD.t46 231.758
R4761 VDD.n361 VDD.n359 206.48
R4762 VDD.n340 VDD.n339 205.865
R4763 VDD.n365 VDD.n364 205.865
R4764 VDD.n363 VDD.n362 205.865
R4765 VDD.n361 VDD.n360 205.865
R4766 VDD.n9 VDD.n8 205.865
R4767 VDD.n7 VDD.n6 205.865
R4768 VDD.n5 VDD.n4 205.865
R4769 VDD.n3 VDD.n2 205.865
R4770 VDD.n28 VDD.n27 205.865
R4771 VDD.n367 VDD.n366 203.143
R4772 VDD.n45 VDD.n44 203.127
R4773 VDD.n26 VDD.n25 203.127
R4774 VDD.n357 VDD.n356 203.127
R4775 VDD.n338 VDD.n337 203.127
R4776 VDD.n43 VDD.n29 203.126
R4777 VDD.n24 VDD.n10 203.126
R4778 VDD.n355 VDD.n341 203.126
R4779 VDD.n336 VDD.n322 203.126
R4780 VDD.n42 VDD.n30 203.03
R4781 VDD.n41 VDD.n40 203.03
R4782 VDD.n23 VDD.n22 203.03
R4783 VDD.n15 VDD.n14 203.03
R4784 VDD.n354 VDD.n342 203.03
R4785 VDD.n353 VDD.n352 203.03
R4786 VDD.n335 VDD.n334 203.03
R4787 VDD.n327 VDD.n326 203.03
R4788 VDD.n189 VDD.n113 185
R4789 VDD.n115 VDD.n113 185
R4790 VDD.n191 VDD.n190 185
R4791 VDD.n192 VDD.n191 185
R4792 VDD.n108 VDD.n107 185
R4793 VDD.n112 VDD.n108 185
R4794 VDD.n201 VDD.n200 185
R4795 VDD.n200 VDD.n199 185
R4796 VDD.n202 VDD.n106 185
R4797 VDD.n198 VDD.n106 185
R4798 VDD.n204 VDD.n203 185
R4799 VDD.n205 VDD.n204 185
R4800 VDD.n101 VDD.n100 185
R4801 VDD.n105 VDD.n101 185
R4802 VDD.n214 VDD.n213 185
R4803 VDD.n213 VDD.n212 185
R4804 VDD.n215 VDD.n99 185
R4805 VDD.n211 VDD.n99 185
R4806 VDD.n217 VDD.n216 185
R4807 VDD.n218 VDD.n217 185
R4808 VDD.n94 VDD.n93 185
R4809 VDD.n98 VDD.n94 185
R4810 VDD.n226 VDD.n225 185
R4811 VDD.n225 VDD.n224 185
R4812 VDD.n227 VDD.n92 185
R4813 VDD.n92 VDD.n91 185
R4814 VDD.n229 VDD.n228 185
R4815 VDD.n230 VDD.n229 185
R4816 VDD.n86 VDD.n85 185
R4817 VDD.n87 VDD.n86 185
R4818 VDD.n238 VDD.n237 185
R4819 VDD.n237 VDD.n236 185
R4820 VDD.n239 VDD.n84 185
R4821 VDD.n84 VDD.n83 185
R4822 VDD.n241 VDD.n240 185
R4823 VDD.n242 VDD.n241 185
R4824 VDD.n78 VDD.n77 185
R4825 VDD.n79 VDD.n78 185
R4826 VDD.n250 VDD.n249 185
R4827 VDD.n249 VDD.n248 185
R4828 VDD.n251 VDD.n76 185
R4829 VDD.n76 VDD.n75 185
R4830 VDD.n253 VDD.n252 185
R4831 VDD.n254 VDD.n253 185
R4832 VDD.n69 VDD.n68 185
R4833 VDD.n70 VDD.n69 185
R4834 VDD.n296 VDD.n295 185
R4835 VDD.n295 VDD.n294 185
R4836 VDD.n297 VDD.n67 185
R4837 VDD.n67 VDD.n53 185
R4838 VDD.n140 VDD.n139 185
R4839 VDD.n141 VDD.n137 185
R4840 VDD.n143 VDD.n142 185
R4841 VDD.n145 VDD.n136 185
R4842 VDD.n147 VDD.n146 185
R4843 VDD.n133 VDD.n132 185
R4844 VDD.n152 VDD.n151 185
R4845 VDD.n154 VDD.n130 185
R4846 VDD.n156 VDD.n155 185
R4847 VDD.n157 VDD.n129 185
R4848 VDD.n159 VDD.n158 185
R4849 VDD.n161 VDD.n127 185
R4850 VDD.n163 VDD.n162 185
R4851 VDD.n164 VDD.n126 185
R4852 VDD.n166 VDD.n165 185
R4853 VDD.n168 VDD.n124 185
R4854 VDD.n170 VDD.n169 185
R4855 VDD.n123 VDD.n121 185
R4856 VDD.n175 VDD.n174 185
R4857 VDD.n177 VDD.n119 185
R4858 VDD.n179 VDD.n178 185
R4859 VDD.n180 VDD.n118 185
R4860 VDD.n182 VDD.n181 185
R4861 VDD.n184 VDD.n117 185
R4862 VDD.n185 VDD.n114 185
R4863 VDD.n188 VDD.n187 185
R4864 VDD.n291 VDD.n72 185
R4865 VDD.n72 VDD.n53 185
R4866 VDD.n293 VDD.n292 185
R4867 VDD.n294 VDD.n293 185
R4868 VDD.n257 VDD.n71 185
R4869 VDD.n71 VDD.n70 185
R4870 VDD.n256 VDD.n255 185
R4871 VDD.n255 VDD.n254 185
R4872 VDD.n74 VDD.n73 185
R4873 VDD.n75 VDD.n74 185
R4874 VDD.n247 VDD.n246 185
R4875 VDD.n248 VDD.n247 185
R4876 VDD.n245 VDD.n80 185
R4877 VDD.n80 VDD.n79 185
R4878 VDD.n244 VDD.n243 185
R4879 VDD.n243 VDD.n242 185
R4880 VDD.n82 VDD.n81 185
R4881 VDD.n83 VDD.n82 185
R4882 VDD.n235 VDD.n234 185
R4883 VDD.n236 VDD.n235 185
R4884 VDD.n233 VDD.n88 185
R4885 VDD.n88 VDD.n87 185
R4886 VDD.n232 VDD.n231 185
R4887 VDD.n231 VDD.n230 185
R4888 VDD.n90 VDD.n89 185
R4889 VDD.n91 VDD.n90 185
R4890 VDD.n223 VDD.n222 185
R4891 VDD.n224 VDD.n223 185
R4892 VDD.n221 VDD.n95 185
R4893 VDD.n98 VDD.n95 185
R4894 VDD.n220 VDD.n219 185
R4895 VDD.n219 VDD.n218 185
R4896 VDD.n97 VDD.n96 185
R4897 VDD.n211 VDD.n97 185
R4898 VDD.n210 VDD.n209 185
R4899 VDD.n212 VDD.n210 185
R4900 VDD.n208 VDD.n102 185
R4901 VDD.n105 VDD.n102 185
R4902 VDD.n207 VDD.n206 185
R4903 VDD.n206 VDD.n205 185
R4904 VDD.n104 VDD.n103 185
R4905 VDD.n198 VDD.n104 185
R4906 VDD.n197 VDD.n196 185
R4907 VDD.n199 VDD.n197 185
R4908 VDD.n195 VDD.n109 185
R4909 VDD.n112 VDD.n109 185
R4910 VDD.n194 VDD.n193 185
R4911 VDD.n193 VDD.n192 185
R4912 VDD.n111 VDD.n110 185
R4913 VDD.n115 VDD.n111 185
R4914 VDD.n312 VDD.n311 185
R4915 VDD.n310 VDD.n66 185
R4916 VDD.n298 VDD.n65 185
R4917 VDD.n314 VDD.n65 185
R4918 VDD.n300 VDD.n299 185
R4919 VDD.n306 VDD.n305 185
R4920 VDD.n304 VDD.n303 185
R4921 VDD.n302 VDD.n301 185
R4922 VDD.n52 VDD.n49 185
R4923 VDD.n317 VDD.n316 185
R4924 VDD.n259 VDD.n51 185
R4925 VDD.n261 VDD.n260 185
R4926 VDD.n263 VDD.n262 185
R4927 VDD.n265 VDD.n264 185
R4928 VDD.n267 VDD.n266 185
R4929 VDD.n269 VDD.n268 185
R4930 VDD.n271 VDD.n270 185
R4931 VDD.n273 VDD.n272 185
R4932 VDD.n275 VDD.n274 185
R4933 VDD.n277 VDD.n276 185
R4934 VDD.n279 VDD.n278 185
R4935 VDD.n281 VDD.n280 185
R4936 VDD.n283 VDD.n282 185
R4937 VDD.n285 VDD.n284 185
R4938 VDD.n287 VDD.n286 185
R4939 VDD.n289 VDD.n288 185
R4940 VDD.n290 VDD.n64 185
R4941 VDD.n314 VDD.n64 185
R4942 VDD.n162 VDD.n128 107.683
R4943 VDD.n128 VDD.n126 107.683
R4944 VDD.n1 VDD.n0 101.662
R4945 VDD.n278 VDD.n61 78.9253
R4946 VDD.n176 VDD.n175 78.9253
R4947 VDD.n177 VDD.n176 78.9253
R4948 VDD.n281 VDD.n61 78.9253
R4949 VDD.n189 VDD.n188 77.177
R4950 VDD.n311 VDD.n297 77.177
R4951 VDD.n140 VDD.n110 77.177
R4952 VDD.n291 VDD.n290 77.177
R4953 VDD.n313 VDD.n312 72.7879
R4954 VDD.n299 VDD.n54 72.7879
R4955 VDD.n304 VDD.n55 72.7879
R4956 VDD.n315 VDD.n52 72.7879
R4957 VDD.n56 VDD.n51 72.7879
R4958 VDD.n262 VDD.n57 72.7879
R4959 VDD.n266 VDD.n58 72.7879
R4960 VDD.n270 VDD.n59 72.7879
R4961 VDD.n274 VDD.n60 72.7879
R4962 VDD.n282 VDD.n62 72.7879
R4963 VDD.n286 VDD.n63 72.7879
R4964 VDD.n186 VDD.n185 72.7879
R4965 VDD.n183 VDD.n182 72.7879
R4966 VDD.n178 VDD.n120 72.7879
R4967 VDD.n169 VDD.n125 72.7879
R4968 VDD.n167 VDD.n166 72.7879
R4969 VDD.n160 VDD.n159 72.7879
R4970 VDD.n155 VDD.n131 72.7879
R4971 VDD.n153 VDD.n152 72.7879
R4972 VDD.n146 VDD.n135 72.7879
R4973 VDD.n144 VDD.n143 72.7879
R4974 VDD.n139 VDD.n138 72.7879
R4975 VDD.n138 VDD.n137 72.7879
R4976 VDD.n145 VDD.n144 72.7879
R4977 VDD.n135 VDD.n132 72.7879
R4978 VDD.n154 VDD.n153 72.7879
R4979 VDD.n131 VDD.n129 72.7879
R4980 VDD.n161 VDD.n160 72.7879
R4981 VDD.n168 VDD.n167 72.7879
R4982 VDD.n125 VDD.n121 72.7879
R4983 VDD.n120 VDD.n118 72.7879
R4984 VDD.n184 VDD.n183 72.7879
R4985 VDD.n187 VDD.n186 72.7879
R4986 VDD.n313 VDD.n66 72.7879
R4987 VDD.n305 VDD.n54 72.7879
R4988 VDD.n301 VDD.n55 72.7879
R4989 VDD.n316 VDD.n315 72.7879
R4990 VDD.n261 VDD.n56 72.7879
R4991 VDD.n265 VDD.n57 72.7879
R4992 VDD.n269 VDD.n58 72.7879
R4993 VDD.n273 VDD.n59 72.7879
R4994 VDD.n277 VDD.n60 72.7879
R4995 VDD.n285 VDD.n62 72.7879
R4996 VDD.n288 VDD.n63 72.7879
R4997 VDD.n116 VDD.n115 57.1093
R4998 VDD.n314 VDD.n53 57.1093
R4999 VDD.n138 VDD.n116 56.1076
R5000 VDD.n144 VDD.n116 56.1076
R5001 VDD.n135 VDD.n116 56.1076
R5002 VDD.n153 VDD.n116 56.1076
R5003 VDD.n131 VDD.n116 56.1076
R5004 VDD.n160 VDD.n116 56.1076
R5005 VDD.n167 VDD.n116 56.1076
R5006 VDD.n125 VDD.n116 56.1076
R5007 VDD.n120 VDD.n116 56.1076
R5008 VDD.n183 VDD.n116 56.1076
R5009 VDD.n186 VDD.n116 56.1076
R5010 VDD.n314 VDD.n313 56.1076
R5011 VDD.n314 VDD.n54 56.1076
R5012 VDD.n314 VDD.n55 56.1076
R5013 VDD.n315 VDD.n314 56.1076
R5014 VDD.n314 VDD.n56 56.1076
R5015 VDD.n314 VDD.n57 56.1076
R5016 VDD.n314 VDD.n58 56.1076
R5017 VDD.n314 VDD.n59 56.1076
R5018 VDD.n314 VDD.n60 56.1076
R5019 VDD.n314 VDD.n62 56.1076
R5020 VDD.n314 VDD.n63 56.1076
R5021 VDD.n164 VDD.n163 54.9652
R5022 VDD.n267 VDD.n264 54.9652
R5023 VDD.n176 VDD.n116 53.0388
R5024 VDD.n314 VDD.n61 53.0388
R5025 VDD.n0 VDD.t68 41.0864
R5026 VDD.n128 VDD.n116 38.6605
R5027 VDD.n192 VDD.n112 30.8211
R5028 VDD.n199 VDD.n198 30.8211
R5029 VDD.n205 VDD.n105 30.8211
R5030 VDD.n212 VDD.n211 30.8211
R5031 VDD.n218 VDD.n98 30.8211
R5032 VDD.n224 VDD.n91 30.8211
R5033 VDD.n230 VDD.n91 30.8211
R5034 VDD.n236 VDD.n87 30.8211
R5035 VDD.n242 VDD.n83 30.8211
R5036 VDD.n248 VDD.n79 30.8211
R5037 VDD.n254 VDD.n75 30.8211
R5038 VDD.n294 VDD.n70 30.8211
R5039 VDD.n98 VDD.t2 30.3679
R5040 VDD.t4 VDD.n87 30.3679
R5041 VDD.n211 VDD.t0 29.4614
R5042 VDD.t8 VDD.n83 29.4614
R5043 VDD.n302 VDD.n49 29.3652
R5044 VDD.n280 VDD.n279 29.3652
R5045 VDD.n8 VDD.t65 28.5655
R5046 VDD.n8 VDD.t74 28.5655
R5047 VDD.n6 VDD.t61 28.5655
R5048 VDD.n6 VDD.t58 28.5655
R5049 VDD.n4 VDD.t70 28.5655
R5050 VDD.n4 VDD.t67 28.5655
R5051 VDD.n2 VDD.t63 28.5655
R5052 VDD.n2 VDD.t73 28.5655
R5053 VDD.t34 VDD.n42 28.5655
R5054 VDD.n42 VDD.t37 28.5655
R5055 VDD.t37 VDD.n41 28.5655
R5056 VDD.n41 VDD.t13 28.5655
R5057 VDD.t55 VDD.n43 28.5655
R5058 VDD.n43 VDD.t34 28.5655
R5059 VDD.n44 VDD.t9 28.5655
R5060 VDD.n44 VDD.t55 28.5655
R5061 VDD.n27 VDD.t7 28.5655
R5062 VDD.n27 VDD.t10 28.5655
R5063 VDD.n23 VDD.t17 28.5655
R5064 VDD.t53 VDD.n23 28.5655
R5065 VDD.n14 VDD.t41 28.5655
R5066 VDD.n14 VDD.t17 28.5655
R5067 VDD.n24 VDD.t53 28.5655
R5068 VDD.t31 VDD.n24 28.5655
R5069 VDD.n25 VDD.t31 28.5655
R5070 VDD.n25 VDD.t6 28.5655
R5071 VDD.n356 VDD.t76 28.5655
R5072 VDD.n356 VDD.t20 28.5655
R5073 VDD.t43 VDD.n354 28.5655
R5074 VDD.n354 VDD.t48 28.5655
R5075 VDD.t48 VDD.n353 28.5655
R5076 VDD.n353 VDD.t25 28.5655
R5077 VDD.t20 VDD.n355 28.5655
R5078 VDD.n355 VDD.t43 28.5655
R5079 VDD.n337 VDD.t39 28.5655
R5080 VDD.n337 VDD.t1 28.5655
R5081 VDD.n335 VDD.t28 28.5655
R5082 VDD.t57 VDD.n335 28.5655
R5083 VDD.n326 VDD.t50 28.5655
R5084 VDD.n326 VDD.t28 28.5655
R5085 VDD.n336 VDD.t57 28.5655
R5086 VDD.t39 VDD.n336 28.5655
R5087 VDD.n339 VDD.t3 28.5655
R5088 VDD.n339 VDD.t5 28.5655
R5089 VDD.n366 VDD.t59 28.5655
R5090 VDD.n366 VDD.t45 28.5655
R5091 VDD.n364 VDD.t64 28.5655
R5092 VDD.n364 VDD.t72 28.5655
R5093 VDD.n362 VDD.t60 28.5655
R5094 VDD.n362 VDD.t75 28.5655
R5095 VDD.n360 VDD.t69 28.5655
R5096 VDD.n360 VDD.t66 28.5655
R5097 VDD.n359 VDD.t62 28.5655
R5098 VDD.n359 VDD.t71 28.5655
R5099 VDD.n105 VDD.t30 28.5549
R5100 VDD.t19 VDD.n79 28.5549
R5101 VDD.n198 VDD.t52 27.6484
R5102 VDD.t33 VDD.n75 27.6484
R5103 VDD.n112 VDD.t16 26.7419
R5104 VDD.t36 VDD.n70 26.7419
R5105 VDD.n115 VDD.t22 25.8354
R5106 VDD.t12 VDD.n53 25.8354
R5107 VDD.n190 VDD.n189 25.6005
R5108 VDD.n190 VDD.n107 25.6005
R5109 VDD.n201 VDD.n107 25.6005
R5110 VDD.n202 VDD.n201 25.6005
R5111 VDD.n203 VDD.n202 25.6005
R5112 VDD.n203 VDD.n100 25.6005
R5113 VDD.n214 VDD.n100 25.6005
R5114 VDD.n215 VDD.n214 25.6005
R5115 VDD.n216 VDD.n215 25.6005
R5116 VDD.n216 VDD.n93 25.6005
R5117 VDD.n226 VDD.n93 25.6005
R5118 VDD.n227 VDD.n226 25.6005
R5119 VDD.n228 VDD.n227 25.6005
R5120 VDD.n228 VDD.n85 25.6005
R5121 VDD.n238 VDD.n85 25.6005
R5122 VDD.n239 VDD.n238 25.6005
R5123 VDD.n240 VDD.n239 25.6005
R5124 VDD.n240 VDD.n77 25.6005
R5125 VDD.n250 VDD.n77 25.6005
R5126 VDD.n251 VDD.n250 25.6005
R5127 VDD.n252 VDD.n251 25.6005
R5128 VDD.n252 VDD.n68 25.6005
R5129 VDD.n296 VDD.n68 25.6005
R5130 VDD.n297 VDD.n296 25.6005
R5131 VDD.n188 VDD.n114 25.6005
R5132 VDD.n117 VDD.n114 25.6005
R5133 VDD.n181 VDD.n117 25.6005
R5134 VDD.n181 VDD.n180 25.6005
R5135 VDD.n180 VDD.n179 25.6005
R5136 VDD.n179 VDD.n119 25.6005
R5137 VDD.n170 VDD.n124 25.6005
R5138 VDD.n165 VDD.n124 25.6005
R5139 VDD.n165 VDD.n164 25.6005
R5140 VDD.n163 VDD.n127 25.6005
R5141 VDD.n158 VDD.n127 25.6005
R5142 VDD.n158 VDD.n157 25.6005
R5143 VDD.n157 VDD.n156 25.6005
R5144 VDD.n156 VDD.n130 25.6005
R5145 VDD.n151 VDD.n130 25.6005
R5146 VDD.n142 VDD.n136 25.6005
R5147 VDD.n142 VDD.n141 25.6005
R5148 VDD.n141 VDD.n140 25.6005
R5149 VDD.n194 VDD.n110 25.6005
R5150 VDD.n195 VDD.n194 25.6005
R5151 VDD.n196 VDD.n195 25.6005
R5152 VDD.n196 VDD.n103 25.6005
R5153 VDD.n207 VDD.n103 25.6005
R5154 VDD.n208 VDD.n207 25.6005
R5155 VDD.n209 VDD.n208 25.6005
R5156 VDD.n209 VDD.n96 25.6005
R5157 VDD.n220 VDD.n96 25.6005
R5158 VDD.n221 VDD.n220 25.6005
R5159 VDD.n222 VDD.n221 25.6005
R5160 VDD.n222 VDD.n89 25.6005
R5161 VDD.n232 VDD.n89 25.6005
R5162 VDD.n233 VDD.n232 25.6005
R5163 VDD.n234 VDD.n233 25.6005
R5164 VDD.n234 VDD.n81 25.6005
R5165 VDD.n244 VDD.n81 25.6005
R5166 VDD.n245 VDD.n244 25.6005
R5167 VDD.n246 VDD.n245 25.6005
R5168 VDD.n246 VDD.n73 25.6005
R5169 VDD.n256 VDD.n73 25.6005
R5170 VDD.n257 VDD.n256 25.6005
R5171 VDD.n292 VDD.n257 25.6005
R5172 VDD.n292 VDD.n291 25.6005
R5173 VDD.n311 VDD.n310 25.6005
R5174 VDD.n300 VDD.n298 25.6005
R5175 VDD.n306 VDD.n303 25.6005
R5176 VDD.n303 VDD.n302 25.6005
R5177 VDD.n260 VDD.n259 25.6005
R5178 VDD.n264 VDD.n263 25.6005
R5179 VDD.n268 VDD.n267 25.6005
R5180 VDD.n271 VDD.n268 25.6005
R5181 VDD.n272 VDD.n271 25.6005
R5182 VDD.n275 VDD.n272 25.6005
R5183 VDD.n276 VDD.n275 25.6005
R5184 VDD.n279 VDD.n276 25.6005
R5185 VDD.n283 VDD.n280 25.6005
R5186 VDD.n284 VDD.n283 25.6005
R5187 VDD.n287 VDD.n284 25.6005
R5188 VDD.n289 VDD.n287 25.6005
R5189 VDD.n290 VDD.n289 25.6005
R5190 VDD.n318 VDD.n317 23.3417
R5191 VDD.n174 VDD.n122 21.0829
R5192 VDD.n150 VDD.n133 21.0829
R5193 VDD.n307 VDD.n300 19.577
R5194 VDD.n173 VDD.n123 17.3181
R5195 VDD.n148 VDD.n147 17.3181
R5196 VDD.n259 VDD.n50 17.3181
R5197 VDD.n171 VDD.n170 15.0593
R5198 VDD.n136 VDD.n134 15.0593
R5199 VDD.n260 VDD.n258 14.3064
R5200 VDD.n0 VDD.t23 14.285
R5201 VDD.n310 VDD.n309 13.5534
R5202 VDD.n309 VDD.n298 12.0476
R5203 VDD.n263 VDD.n258 11.2946
R5204 VDD.n171 VDD.n123 10.5417
R5205 VDD.n147 VDD.n134 10.5417
R5206 VDD.n309 VDD.n308 9.43153
R5207 VDD.n258 VDD.n48 9.43153
R5208 VDD.n172 VDD.n122 9.36774
R5209 VDD.n150 VDD.n149 9.36774
R5210 VDD.n172 VDD.n171 9.36429
R5211 VDD.n149 VDD.n134 9.36429
R5212 VDD.n149 VDD.n148 9.3005
R5213 VDD.n173 VDD.n172 9.3005
R5214 VDD.n308 VDD.n307 9.3005
R5215 VDD.n303 VDD.n47 9.3005
R5216 VDD.n319 VDD.n318 9.3005
R5217 VDD.n50 VDD.n48 9.3005
R5218 VDD.n122 VDD.n119 8.28285
R5219 VDD.n174 VDD.n173 8.28285
R5220 VDD.n151 VDD.n150 8.28285
R5221 VDD.n148 VDD.n133 8.28285
R5222 VDD.n317 VDD.n50 8.28285
R5223 VDD.n307 VDD.n306 6.02403
R5224 VDD.n192 VDD.t22 4.98619
R5225 VDD.n294 VDD.t12 4.98619
R5226 VDD.n199 VDD.t16 4.0797
R5227 VDD.n254 VDD.t36 4.0797
R5228 VDD.n28 VDD.n26 3.35217
R5229 VDD.n340 VDD.n338 3.35217
R5230 VDD.n205 VDD.t52 3.17321
R5231 VDD.n248 VDD.t33 3.17321
R5232 VDD.n3 VDD.n1 3.06997
R5233 VDD.n46 VDD.n45 2.73818
R5234 VDD.n358 VDD.n357 2.73818
R5235 VDD.n369 VDD.n368 2.45598
R5236 VDD.n212 VDD.t30 2.26672
R5237 VDD.n242 VDD.t19 2.26672
R5238 VDD.n318 VDD.n49 2.25932
R5239 VDD.n321 VDD.n320 2.20937
R5240 VDD.n370 VDD.n358 2.07758
R5241 VDD.n372 VDD.n9 1.82938
R5242 VDD.n370 VDD.n369 1.63948
R5243 VDD VDD.n372 1.52224
R5244 VDD.n321 VDD.n46 1.485
R5245 VDD.n218 VDD.t0 1.36023
R5246 VDD.n236 VDD.t8 1.36023
R5247 VDD.n371 VDD.n370 0.9725
R5248 VDD.n5 VDD.n3 0.61449
R5249 VDD.n7 VDD.n5 0.61449
R5250 VDD.n9 VDD.n7 0.61449
R5251 VDD.n46 VDD.n28 0.61449
R5252 VDD.n358 VDD.n340 0.61449
R5253 VDD.n363 VDD.n361 0.61449
R5254 VDD.n365 VDD.n363 0.61449
R5255 VDD.n369 VDD.n365 0.61449
R5256 VDD.n371 VDD.n321 0.590949
R5257 VDD.n372 VDD.n371 0.4545
R5258 VDD.n224 VDD.t2 0.453744
R5259 VDD.n230 VDD.t4 0.453744
R5260 VDD.n352 VDD.n343 0.38373
R5261 VDD.n347 VDD.n342 0.38373
R5262 VDD.n328 VDD.n327 0.38373
R5263 VDD.n334 VDD.n323 0.38373
R5264 VDD.n40 VDD.n39 0.383729
R5265 VDD.n33 VDD.n30 0.383729
R5266 VDD.n15 VDD.n13 0.383729
R5267 VDD.n22 VDD.n21 0.383729
R5268 VDD.n35 VDD.n31 0.338735
R5269 VDD.n35 VDD.n29 0.338735
R5270 VDD.n45 VDD.n29 0.338735
R5271 VDD.n16 VDD.n11 0.338735
R5272 VDD.n11 VDD.n10 0.338735
R5273 VDD.n26 VDD.n10 0.338735
R5274 VDD.n351 VDD.n344 0.338735
R5275 VDD.n344 VDD.n341 0.338735
R5276 VDD.n357 VDD.n341 0.338735
R5277 VDD.n333 VDD.n324 0.338735
R5278 VDD.n333 VDD.n322 0.338735
R5279 VDD.n338 VDD.n322 0.338735
R5280 VDD.n38 VDD.n31 0.285826
R5281 VDD.n36 VDD.n35 0.285826
R5282 VDD.n17 VDD.n16 0.285826
R5283 VDD.n19 VDD.n11 0.285826
R5284 VDD.n351 VDD.n350 0.285826
R5285 VDD.n345 VDD.n344 0.285826
R5286 VDD.n325 VDD.n324 0.285826
R5287 VDD.n333 VDD.n332 0.285826
R5288 VDD.n37 VDD.n36 0.188
R5289 VDD.n38 VDD.n37 0.188
R5290 VDD.n34 VDD.n33 0.188
R5291 VDD.n33 VDD.n32 0.188
R5292 VDD.n39 VDD.n32 0.188
R5293 VDD.n18 VDD.n17 0.188
R5294 VDD.n19 VDD.n18 0.188
R5295 VDD.n13 VDD.n12 0.188
R5296 VDD.n21 VDD.n12 0.188
R5297 VDD.n21 VDD.n20 0.188
R5298 VDD.n347 VDD.n346 0.188
R5299 VDD.n348 VDD.n347 0.188
R5300 VDD.n348 VDD.n343 0.188
R5301 VDD.n349 VDD.n345 0.188
R5302 VDD.n350 VDD.n349 0.188
R5303 VDD.n329 VDD.n328 0.188
R5304 VDD.n329 VDD.n323 0.188
R5305 VDD.n331 VDD.n323 0.188
R5306 VDD.n330 VDD.n325 0.188
R5307 VDD.n332 VDD.n330 0.188
R5308 VDD.n40 VDD.n31 0.0984044
R5309 VDD.n35 VDD.n30 0.0984044
R5310 VDD.n16 VDD.n15 0.0984044
R5311 VDD.n22 VDD.n11 0.0984044
R5312 VDD.n344 VDD.n342 0.0984028
R5313 VDD.n352 VDD.n351 0.0984028
R5314 VDD.n334 VDD.n333 0.0984028
R5315 VDD.n327 VDD.n324 0.0984028
R5316 VDD.n368 VDD.n367 0.0793043
R5317 VDD.n308 VDD.n47 0.0729138
R5318 VDD.n319 VDD.n48 0.0729138
R5319 VDD.n320 VDD.n319 0.0686034
R5320 VDD.n320 VDD.n47 0.063431
R5321 a_2080_2896.n87 a_2080_2896.n86 185
R5322 a_2080_2896.n86 a_2080_2896.n85 185
R5323 a_2080_2896.n86 a_2080_2896.n8 185
R5324 a_2080_2896.n86 a_2080_2896.n7 185
R5325 a_2080_2896.n86 a_2080_2896.n6 185
R5326 a_2080_2896.n86 a_2080_2896.n5 185
R5327 a_2080_2896.n86 a_2080_2896.n4 185
R5328 a_2080_2896.n53 a_2080_2896.n52 185
R5329 a_2080_2896.n53 a_2080_2896.n40 185
R5330 a_2080_2896.n53 a_2080_2896.n39 185
R5331 a_2080_2896.n53 a_2080_2896.n37 185
R5332 a_2080_2896.n53 a_2080_2896.n36 185
R5333 a_2080_2896.n54 a_2080_2896.n53 185
R5334 a_2080_2896.t2 a_2080_2896.n92 180.167
R5335 a_2080_2896.t2 a_2080_2896.n92 180.167
R5336 a_2080_2896.n21 a_2080_2896.t35 165.607
R5337 a_2080_2896.n9 a_2080_2896.t22 165.607
R5338 a_2080_2896.n70 a_2080_2896.t20 165.032
R5339 a_2080_2896.n19 a_2080_2896.t21 165.032
R5340 a_2080_2896.n18 a_2080_2896.t8 165.032
R5341 a_2080_2896.n17 a_2080_2896.t18 165.032
R5342 a_2080_2896.n16 a_2080_2896.t29 165.032
R5343 a_2080_2896.n15 a_2080_2896.t28 165.032
R5344 a_2080_2896.n14 a_2080_2896.t39 165.032
R5345 a_2080_2896.n13 a_2080_2896.t40 165.032
R5346 a_2080_2896.n12 a_2080_2896.t11 165.032
R5347 a_2080_2896.n11 a_2080_2896.t10 165.032
R5348 a_2080_2896.n10 a_2080_2896.t9 165.032
R5349 a_2080_2896.n9 a_2080_2896.t30 165.032
R5350 a_2080_2896.n68 a_2080_2896.t42 163.058
R5351 a_2080_2896.n66 a_2080_2896.t31 163.058
R5352 a_2080_2896.n64 a_2080_2896.t41 163.058
R5353 a_2080_2896.n62 a_2080_2896.t13 163.058
R5354 a_2080_2896.n60 a_2080_2896.t12 163.058
R5355 a_2080_2896.n32 a_2080_2896.t25 163.058
R5356 a_2080_2896.n58 a_2080_2896.t23 163.058
R5357 a_2080_2896.n28 a_2080_2896.t34 163.058
R5358 a_2080_2896.n26 a_2080_2896.t33 163.058
R5359 a_2080_2896.n24 a_2080_2896.t32 163.058
R5360 a_2080_2896.n22 a_2080_2896.t15 163.058
R5361 a_2080_2896.n20 a_2080_2896.t43 163.058
R5362 a_2080_2896.t3 a_2080_2896.n56 162.941
R5363 a_2080_2896.n56 a_2080_2896.t5 162.941
R5364 a_2080_2896.n68 a_2080_2896.t26 162.781
R5365 a_2080_2896.n66 a_2080_2896.t14 162.781
R5366 a_2080_2896.n64 a_2080_2896.t24 162.781
R5367 a_2080_2896.n62 a_2080_2896.t37 162.781
R5368 a_2080_2896.n60 a_2080_2896.t36 162.781
R5369 a_2080_2896.n28 a_2080_2896.t19 162.781
R5370 a_2080_2896.n26 a_2080_2896.t17 162.781
R5371 a_2080_2896.n24 a_2080_2896.t16 162.781
R5372 a_2080_2896.n22 a_2080_2896.t38 162.781
R5373 a_2080_2896.n20 a_2080_2896.t27 162.781
R5374 a_2080_2896.n57 a_2080_2896.t3 162.639
R5375 a_2080_2896.t5 a_2080_2896.n33 162.639
R5376 a_2080_2896.n91 a_2080_2896.t0 130.75
R5377 a_2080_2896.n86 a_2080_2896.n3 86.5152
R5378 a_2080_2896.n53 a_2080_2896.n38 86.5152
R5379 a_2080_2896.n88 a_2080_2896.n0 30.3012
R5380 a_2080_2896.n73 a_2080_2896.n4 24.8476
R5381 a_2080_2896.n46 a_2080_2896.n39 24.8476
R5382 a_2080_2896.n44 a_2080_2896.n37 24.8476
R5383 a_2080_2896.n75 a_2080_2896.n5 23.3417
R5384 a_2080_2896.n48 a_2080_2896.n40 23.3417
R5385 a_2080_2896.n42 a_2080_2896.n36 23.3417
R5386 a_2080_2896.n72 a_2080_2896.n3 22.0256
R5387 a_2080_2896.n77 a_2080_2896.n6 21.8358
R5388 a_2080_2896.n52 a_2080_2896.n51 21.8358
R5389 a_2080_2896.n54 a_2080_2896.n35 21.8358
R5390 a_2080_2896.n79 a_2080_2896.n7 20.3299
R5391 a_2080_2896.n81 a_2080_2896.n8 18.824
R5392 a_2080_2896.n85 a_2080_2896.n84 17.3181
R5393 a_2080_2896.n86 a_2080_2896.n0 16.3559
R5394 a_2080_2896.n87 a_2080_2896.n2 15.8123
R5395 a_2080_2896.n52 a_2080_2896.n41 14.5711
R5396 a_2080_2896.n55 a_2080_2896.n54 14.5711
R5397 a_2080_2896.n72 a_2080_2896.n71 12.9589
R5398 a_2080_2896.n73 a_2080_2896.n3 12.7256
R5399 a_2080_2896.n46 a_2080_2896.n38 12.7256
R5400 a_2080_2896.n44 a_2080_2896.n38 12.7256
R5401 a_2080_2896.n88 a_2080_2896.n87 11.2946
R5402 a_2080_2896.n85 a_2080_2896.n2 9.78874
R5403 a_2080_2896.n47 a_2080_2896.n46 9.3005
R5404 a_2080_2896.n49 a_2080_2896.n48 9.3005
R5405 a_2080_2896.n51 a_2080_2896.n50 9.3005
R5406 a_2080_2896.n45 a_2080_2896.n44 9.3005
R5407 a_2080_2896.n43 a_2080_2896.n42 9.3005
R5408 a_2080_2896.n35 a_2080_2896.n34 9.3005
R5409 a_2080_2896.n74 a_2080_2896.n73 9.3005
R5410 a_2080_2896.n76 a_2080_2896.n75 9.3005
R5411 a_2080_2896.n78 a_2080_2896.n77 9.3005
R5412 a_2080_2896.n80 a_2080_2896.n79 9.3005
R5413 a_2080_2896.n82 a_2080_2896.n81 9.3005
R5414 a_2080_2896.n84 a_2080_2896.n83 9.3005
R5415 a_2080_2896.n2 a_2080_2896.n1 9.3005
R5416 a_2080_2896.n89 a_2080_2896.n88 9.3005
R5417 a_2080_2896.n71 a_2080_2896.n70 8.61608
R5418 a_2080_2896.n84 a_2080_2896.n8 8.28285
R5419 a_2080_2896.n81 a_2080_2896.n7 6.77697
R5420 a_2080_2896.n53 a_2080_2896.t6 5.8005
R5421 a_2080_2896.n53 a_2080_2896.t4 5.8005
R5422 a_2080_2896.n79 a_2080_2896.n6 5.27109
R5423 a_2080_2896.n77 a_2080_2896.n5 3.76521
R5424 a_2080_2896.n51 a_2080_2896.n40 3.76521
R5425 a_2080_2896.n36 a_2080_2896.n35 3.76521
R5426 a_2080_2896.n86 a_2080_2896.t7 2.48621
R5427 a_2080_2896.n86 a_2080_2896.t1 2.48621
R5428 a_2080_2896.n90 a_2080_2896.n0 2.36936
R5429 a_2080_2896.n75 a_2080_2896.n4 2.25932
R5430 a_2080_2896.n48 a_2080_2896.n39 2.25932
R5431 a_2080_2896.n42 a_2080_2896.n37 2.25932
R5432 a_2080_2896.n69 a_2080_2896.n68 2.25162
R5433 a_2080_2896.n67 a_2080_2896.n66 2.25162
R5434 a_2080_2896.n65 a_2080_2896.n64 2.25162
R5435 a_2080_2896.n63 a_2080_2896.n62 2.25162
R5436 a_2080_2896.n61 a_2080_2896.n60 2.25162
R5437 a_2080_2896.n32 a_2080_2896.n30 2.25162
R5438 a_2080_2896.n59 a_2080_2896.n58 2.25162
R5439 a_2080_2896.n29 a_2080_2896.n28 2.25162
R5440 a_2080_2896.n27 a_2080_2896.n26 2.25162
R5441 a_2080_2896.n25 a_2080_2896.n24 2.25162
R5442 a_2080_2896.n23 a_2080_2896.n22 2.25162
R5443 a_2080_2896.n21 a_2080_2896.n20 2.25162
R5444 a_2080_2896.n71 a_2080_2896.n19 2.17137
R5445 a_2080_2896.n92 a_2080_2896.n91 1.27148
R5446 a_2080_2896.n23 a_2080_2896.n21 0.574917
R5447 a_2080_2896.n25 a_2080_2896.n23 0.574917
R5448 a_2080_2896.n27 a_2080_2896.n25 0.574917
R5449 a_2080_2896.n29 a_2080_2896.n27 0.574917
R5450 a_2080_2896.n30 a_2080_2896.n29 0.574917
R5451 a_2080_2896.n59 a_2080_2896.n30 0.574917
R5452 a_2080_2896.n61 a_2080_2896.n59 0.574917
R5453 a_2080_2896.n63 a_2080_2896.n61 0.574917
R5454 a_2080_2896.n65 a_2080_2896.n63 0.574917
R5455 a_2080_2896.n67 a_2080_2896.n65 0.574917
R5456 a_2080_2896.n69 a_2080_2896.n67 0.574917
R5457 a_2080_2896.n70 a_2080_2896.n69 0.574917
R5458 a_2080_2896.n10 a_2080_2896.n9 0.574917
R5459 a_2080_2896.n11 a_2080_2896.n10 0.574917
R5460 a_2080_2896.n12 a_2080_2896.n11 0.574917
R5461 a_2080_2896.n13 a_2080_2896.n12 0.574917
R5462 a_2080_2896.n14 a_2080_2896.n13 0.574917
R5463 a_2080_2896.n15 a_2080_2896.n14 0.574917
R5464 a_2080_2896.n16 a_2080_2896.n15 0.574917
R5465 a_2080_2896.n17 a_2080_2896.n16 0.574917
R5466 a_2080_2896.n18 a_2080_2896.n17 0.574917
R5467 a_2080_2896.n19 a_2080_2896.n18 0.574917
R5468 a_2080_2896.n91 a_2080_2896.n90 0.320353
R5469 a_2080_2896.n33 a_2080_2896.n31 0.302413
R5470 a_2080_2896.n57 a_2080_2896.n31 0.302413
R5471 a_2080_2896.n41 a_2080_2896.n31 0.217891
R5472 a_2080_2896.n56 a_2080_2896.n55 0.217891
R5473 a_2080_2896.n50 a_2080_2896.n41 0.196152
R5474 a_2080_2896.n50 a_2080_2896.n49 0.196152
R5475 a_2080_2896.n49 a_2080_2896.n47 0.196152
R5476 a_2080_2896.n47 a_2080_2896.n45 0.196152
R5477 a_2080_2896.n45 a_2080_2896.n43 0.196152
R5478 a_2080_2896.n43 a_2080_2896.n34 0.196152
R5479 a_2080_2896.n55 a_2080_2896.n34 0.196152
R5480 a_2080_2896.n90 a_2080_2896.n89 0.196152
R5481 a_2080_2896.n89 a_2080_2896.n1 0.196152
R5482 a_2080_2896.n83 a_2080_2896.n1 0.196152
R5483 a_2080_2896.n83 a_2080_2896.n82 0.196152
R5484 a_2080_2896.n82 a_2080_2896.n80 0.196152
R5485 a_2080_2896.n80 a_2080_2896.n78 0.196152
R5486 a_2080_2896.n78 a_2080_2896.n76 0.196152
R5487 a_2080_2896.n76 a_2080_2896.n74 0.196152
R5488 a_2080_2896.n74 a_2080_2896.n72 0.196152
R5489 a_2080_2896.n33 a_2080_2896.n32 0.142018
R5490 a_2080_2896.n58 a_2080_2896.n57 0.142018
R5491 a_4920_2896.n46 a_4920_2896.n28 185
R5492 a_4920_2896.n46 a_4920_2896.n27 185
R5493 a_4920_2896.n46 a_4920_2896.n26 185
R5494 a_4920_2896.n46 a_4920_2896.n25 185
R5495 a_4920_2896.n46 a_4920_2896.n24 185
R5496 a_4920_2896.n46 a_4920_2896.n23 185
R5497 a_4920_2896.n46 a_4920_2896.n22 185
R5498 a_4920_2896.n30 a_4920_2896.t25 130.75
R5499 a_4920_2896.n30 a_4920_2896.t26 91.3557
R5500 a_4920_2896.n47 a_4920_2896.n46 86.5152
R5501 a_4920_2896.n45 a_4920_2896.n29 30.3012
R5502 a_4920_2896.n15 a_4920_2896.n14 26.8581
R5503 a_4920_2896.n5 a_4920_2896.n4 26.6299
R5504 a_4920_2896.n19 a_4920_2896.n9 25.7063
R5505 a_4920_2896.n18 a_4920_2896.n10 25.7063
R5506 a_4920_2896.n17 a_4920_2896.n11 25.7063
R5507 a_4920_2896.n16 a_4920_2896.n12 25.7063
R5508 a_4920_2896.n15 a_4920_2896.n13 25.7063
R5509 a_4920_2896.n51 a_4920_2896.n50 25.4783
R5510 a_4920_2896.n5 a_4920_2896.n3 25.4781
R5511 a_4920_2896.n6 a_4920_2896.n2 25.4781
R5512 a_4920_2896.n7 a_4920_2896.n1 25.4781
R5513 a_4920_2896.n8 a_4920_2896.n0 25.4781
R5514 a_4920_2896.n22 a_4920_2896.n21 24.8476
R5515 a_4920_2896.n31 a_4920_2896.n23 23.3417
R5516 a_4920_2896.n48 a_4920_2896.n47 22.0256
R5517 a_4920_2896.n33 a_4920_2896.n24 21.8358
R5518 a_4920_2896.n35 a_4920_2896.n25 20.3299
R5519 a_4920_2896.n37 a_4920_2896.n26 18.824
R5520 a_4920_2896.n39 a_4920_2896.n27 17.3181
R5521 a_4920_2896.n46 a_4920_2896.n45 16.3559
R5522 a_4920_2896.n41 a_4920_2896.n28 15.8123
R5523 a_4920_2896.n47 a_4920_2896.n21 12.7256
R5524 a_4920_2896.n29 a_4920_2896.n28 11.2946
R5525 a_4920_2896.n41 a_4920_2896.n27 9.78874
R5526 a_4920_2896.n49 a_4920_2896.n19 9.30285
R5527 a_4920_2896.n21 a_4920_2896.n20 9.3005
R5528 a_4920_2896.n32 a_4920_2896.n31 9.3005
R5529 a_4920_2896.n34 a_4920_2896.n33 9.3005
R5530 a_4920_2896.n36 a_4920_2896.n35 9.3005
R5531 a_4920_2896.n38 a_4920_2896.n37 9.3005
R5532 a_4920_2896.n40 a_4920_2896.n39 9.3005
R5533 a_4920_2896.n42 a_4920_2896.n41 9.3005
R5534 a_4920_2896.n43 a_4920_2896.n29 9.3005
R5535 a_4920_2896.n39 a_4920_2896.n26 8.28285
R5536 a_4920_2896.n37 a_4920_2896.n25 6.77697
R5537 a_4920_2896.n4 a_4920_2896.t14 5.8005
R5538 a_4920_2896.n4 a_4920_2896.t9 5.8005
R5539 a_4920_2896.n3 a_4920_2896.t22 5.8005
R5540 a_4920_2896.n3 a_4920_2896.t21 5.8005
R5541 a_4920_2896.n2 a_4920_2896.t20 5.8005
R5542 a_4920_2896.n2 a_4920_2896.t3 5.8005
R5543 a_4920_2896.n1 a_4920_2896.t4 5.8005
R5544 a_4920_2896.n1 a_4920_2896.t11 5.8005
R5545 a_4920_2896.n0 a_4920_2896.t10 5.8005
R5546 a_4920_2896.n0 a_4920_2896.t16 5.8005
R5547 a_4920_2896.n9 a_4920_2896.t8 5.8005
R5548 a_4920_2896.n9 a_4920_2896.t1 5.8005
R5549 a_4920_2896.n10 a_4920_2896.t18 5.8005
R5550 a_4920_2896.n10 a_4920_2896.t2 5.8005
R5551 a_4920_2896.n11 a_4920_2896.t13 5.8005
R5552 a_4920_2896.n11 a_4920_2896.t19 5.8005
R5553 a_4920_2896.n12 a_4920_2896.t5 5.8005
R5554 a_4920_2896.n12 a_4920_2896.t12 5.8005
R5555 a_4920_2896.n13 a_4920_2896.t7 5.8005
R5556 a_4920_2896.n13 a_4920_2896.t6 5.8005
R5557 a_4920_2896.n14 a_4920_2896.t0 5.8005
R5558 a_4920_2896.n14 a_4920_2896.t17 5.8005
R5559 a_4920_2896.t23 a_4920_2896.n51 5.8005
R5560 a_4920_2896.n51 a_4920_2896.t15 5.8005
R5561 a_4920_2896.n35 a_4920_2896.n24 5.27109
R5562 a_4920_2896.n33 a_4920_2896.n23 3.76521
R5563 a_4920_2896.n50 a_4920_2896.n49 2.92217
R5564 a_4920_2896.n46 a_4920_2896.t26 2.48621
R5565 a_4920_2896.n46 a_4920_2896.t24 2.48621
R5566 a_4920_2896.n45 a_4920_2896.n44 2.36936
R5567 a_4920_2896.n31 a_4920_2896.n22 2.25932
R5568 a_4920_2896.n49 a_4920_2896.n48 2.19829
R5569 a_4920_2896.n16 a_4920_2896.n15 1.15229
R5570 a_4920_2896.n17 a_4920_2896.n16 1.15229
R5571 a_4920_2896.n18 a_4920_2896.n17 1.15229
R5572 a_4920_2896.n19 a_4920_2896.n18 1.15229
R5573 a_4920_2896.n6 a_4920_2896.n5 1.15229
R5574 a_4920_2896.n7 a_4920_2896.n6 1.15229
R5575 a_4920_2896.n8 a_4920_2896.n7 1.15229
R5576 a_4920_2896.n50 a_4920_2896.n8 1.15229
R5577 a_4920_2896.n44 a_4920_2896.n30 0.320353
R5578 a_4920_2896.n44 a_4920_2896.n43 0.196152
R5579 a_4920_2896.n43 a_4920_2896.n42 0.196152
R5580 a_4920_2896.n42 a_4920_2896.n40 0.196152
R5581 a_4920_2896.n40 a_4920_2896.n38 0.196152
R5582 a_4920_2896.n38 a_4920_2896.n36 0.196152
R5583 a_4920_2896.n36 a_4920_2896.n34 0.196152
R5584 a_4920_2896.n34 a_4920_2896.n32 0.196152
R5585 a_4920_2896.n32 a_4920_2896.n20 0.196152
R5586 a_4920_2896.n48 a_4920_2896.n20 0.196152
R5587 VP.n0 VP.t7 263.647
R5588 VP.n3 VP.t3 262.863
R5589 VP.n2 VP.t1 262.498
R5590 VP.n0 VP.t6 261.709
R5591 VP.n1 VP.t2 261.709
R5592 VP.n3 VP.t5 261.584
R5593 VP.n4 VP.t4 261.584
R5594 VP.n5 VP.t0 261.433
R5595 VP.n6 VP.n2 8.91083
R5596 VP VP.n6 2.38312
R5597 VP.n1 VP.n0 1.72698
R5598 VP.n6 VP.n5 1.52193
R5599 VP.n5 VP.n4 1.4312
R5600 VP.n4 VP.n3 1.16675
R5601 VP.n2 VP.n1 1.14999
R5602 a_2995_7336.n30 a_2995_7336.n29 185
R5603 a_2995_7336.n30 a_2995_7336.n12 185
R5604 a_2995_7336.n30 a_2995_7336.n11 185
R5605 a_2995_7336.n30 a_2995_7336.n10 185
R5606 a_2995_7336.n30 a_2995_7336.n9 185
R5607 a_2995_7336.n30 a_2995_7336.n8 185
R5608 a_2995_7336.n30 a_2995_7336.n7 185
R5609 a_2995_7336.n13 a_2995_7336.t5 130.75
R5610 a_2995_7336.n13 a_2995_7336.t7 91.3557
R5611 a_2995_7336.n31 a_2995_7336.n30 86.5152
R5612 a_2995_7336.n15 a_2995_7336.n6 30.3012
R5613 a_2995_7336.n29 a_2995_7336.n5 24.8476
R5614 a_2995_7336.n28 a_2995_7336.n12 23.3417
R5615 a_2995_7336.n32 a_2995_7336.n31 22.0256
R5616 a_2995_7336.n25 a_2995_7336.n11 21.8358
R5617 a_2995_7336.n23 a_2995_7336.n10 20.3299
R5618 a_2995_7336.n21 a_2995_7336.n9 18.824
R5619 a_2995_7336.n19 a_2995_7336.n8 17.3181
R5620 a_2995_7336.n30 a_2995_7336.n6 16.3559
R5621 a_2995_7336.n17 a_2995_7336.n7 15.8123
R5622 a_2995_7336.n31 a_2995_7336.n5 12.7256
R5623 a_2995_7336.n39 a_2995_7336.n38 12.1709
R5624 a_2995_7336.n40 a_2995_7336.n39 12.1709
R5625 a_2995_7336.n40 a_2995_7336.n0 11.493
R5626 a_2995_7336.n38 a_2995_7336.n33 11.493
R5627 a_2995_7336.n37 a_2995_7336.n35 11.493
R5628 a_2995_7336.n3 a_2995_7336.n1 11.493
R5629 a_2995_7336.n41 a_2995_7336.n40 11.493
R5630 a_2995_7336.n38 a_2995_7336.n34 11.4929
R5631 a_2995_7336.n37 a_2995_7336.n36 11.4929
R5632 a_2995_7336.n3 a_2995_7336.n2 11.4929
R5633 a_2995_7336.n15 a_2995_7336.n7 11.2946
R5634 a_2995_7336.n17 a_2995_7336.n8 9.78874
R5635 a_2995_7336.n5 a_2995_7336.n4 9.3005
R5636 a_2995_7336.n28 a_2995_7336.n27 9.3005
R5637 a_2995_7336.n26 a_2995_7336.n25 9.3005
R5638 a_2995_7336.n24 a_2995_7336.n23 9.3005
R5639 a_2995_7336.n22 a_2995_7336.n21 9.3005
R5640 a_2995_7336.n20 a_2995_7336.n19 9.3005
R5641 a_2995_7336.n18 a_2995_7336.n17 9.3005
R5642 a_2995_7336.n16 a_2995_7336.n15 9.3005
R5643 a_2995_7336.n19 a_2995_7336.n9 8.28285
R5644 a_2995_7336.n21 a_2995_7336.n10 6.77697
R5645 a_2995_7336.n23 a_2995_7336.n11 5.27109
R5646 a_2995_7336.n25 a_2995_7336.n12 3.76521
R5647 a_2995_7336.n39 a_2995_7336.n32 3.48602
R5648 a_2995_7336.n0 a_2995_7336.t10 2.48621
R5649 a_2995_7336.n0 a_2995_7336.t1 2.48621
R5650 a_2995_7336.n34 a_2995_7336.t17 2.48621
R5651 a_2995_7336.n34 a_2995_7336.t9 2.48621
R5652 a_2995_7336.n33 a_2995_7336.t19 2.48621
R5653 a_2995_7336.n33 a_2995_7336.t16 2.48621
R5654 a_2995_7336.n36 a_2995_7336.t8 2.48621
R5655 a_2995_7336.n36 a_2995_7336.t13 2.48621
R5656 a_2995_7336.n35 a_2995_7336.t15 2.48621
R5657 a_2995_7336.n35 a_2995_7336.t3 2.48621
R5658 a_2995_7336.n2 a_2995_7336.t12 2.48621
R5659 a_2995_7336.n2 a_2995_7336.t4 2.48621
R5660 a_2995_7336.n1 a_2995_7336.t18 2.48621
R5661 a_2995_7336.n1 a_2995_7336.t11 2.48621
R5662 a_2995_7336.n30 a_2995_7336.t2 2.48621
R5663 a_2995_7336.n30 a_2995_7336.t6 2.48621
R5664 a_2995_7336.t0 a_2995_7336.n41 2.48621
R5665 a_2995_7336.n41 a_2995_7336.t14 2.48621
R5666 a_2995_7336.n14 a_2995_7336.n6 2.36936
R5667 a_2995_7336.n29 a_2995_7336.n28 2.25932
R5668 a_2995_7336.n38 a_2995_7336.n37 1.15229
R5669 a_2995_7336.n37 a_2995_7336.n3 1.15229
R5670 a_2995_7336.n40 a_2995_7336.n3 1.15229
R5671 a_2995_7336.n14 a_2995_7336.n13 0.320353
R5672 a_2995_7336.n32 a_2995_7336.n4 0.196152
R5673 a_2995_7336.n27 a_2995_7336.n4 0.196152
R5674 a_2995_7336.n27 a_2995_7336.n26 0.196152
R5675 a_2995_7336.n26 a_2995_7336.n24 0.196152
R5676 a_2995_7336.n24 a_2995_7336.n22 0.196152
R5677 a_2995_7336.n22 a_2995_7336.n20 0.196152
R5678 a_2995_7336.n20 a_2995_7336.n18 0.196152
R5679 a_2995_7336.n18 a_2995_7336.n16 0.196152
R5680 a_2995_7336.n16 a_2995_7336.n14 0.196152
R5681 VN.n0 VN.t0 263.647
R5682 VN.n3 VN.t2 262.863
R5683 VN.n2 VN.t5 262.498
R5684 VN.n1 VN.t4 261.709
R5685 VN.n0 VN.t1 261.709
R5686 VN.n4 VN.t7 261.584
R5687 VN.n3 VN.t6 261.584
R5688 VN.n5 VN.t3 261.433
R5689 VN.n6 VN.n2 8.91083
R5690 VN VN.n6 2.48729
R5691 VN.n1 VN.n0 1.72698
R5692 VN.n6 VN.n5 1.52193
R5693 VN.n5 VN.n4 1.4312
R5694 VN.n4 VN.n3 1.16675
R5695 VN.n2 VN.n1 1.14999
R5696 a_2479_9004.n70 a_2479_9004.t22 260.111
R5697 a_2479_9004.n4 a_2479_9004.t21 260.111
R5698 a_2479_9004.n3 a_2479_9004.t0 260.111
R5699 a_2479_9004.n1 a_2479_9004.t2 260.111
R5700 a_2479_9004.n70 a_2479_9004.t4 260.111
R5701 a_2479_9004.n4 a_2479_9004.t6 260.111
R5702 a_2479_9004.n3 a_2479_9004.t24 260.111
R5703 a_2479_9004.n1 a_2479_9004.t23 260.111
R5704 a_2479_9004.n2 a_2479_9004.n0 203.413
R5705 a_2479_9004.n72 a_2479_9004.n71 203.412
R5706 a_2479_9004.n34 a_2479_9004.n33 185
R5707 a_2479_9004.n34 a_2479_9004.n16 185
R5708 a_2479_9004.n34 a_2479_9004.n15 185
R5709 a_2479_9004.n34 a_2479_9004.n14 185
R5710 a_2479_9004.n34 a_2479_9004.n13 185
R5711 a_2479_9004.n34 a_2479_9004.n12 185
R5712 a_2479_9004.n34 a_2479_9004.n11 185
R5713 a_2479_9004.n65 a_2479_9004.n64 185
R5714 a_2479_9004.n65 a_2479_9004.n47 185
R5715 a_2479_9004.n65 a_2479_9004.n46 185
R5716 a_2479_9004.n65 a_2479_9004.n45 185
R5717 a_2479_9004.n65 a_2479_9004.n44 185
R5718 a_2479_9004.n65 a_2479_9004.n43 185
R5719 a_2479_9004.n65 a_2479_9004.n42 185
R5720 a_2479_9004.n17 a_2479_9004.t8 130.75
R5721 a_2479_9004.n48 a_2479_9004.t11 130.75
R5722 a_2479_9004.n17 a_2479_9004.t10 91.3557
R5723 a_2479_9004.n48 a_2479_9004.t12 91.3557
R5724 a_2479_9004.n35 a_2479_9004.n34 86.5152
R5725 a_2479_9004.n66 a_2479_9004.n65 86.5152
R5726 a_2479_9004.n19 a_2479_9004.n10 30.3012
R5727 a_2479_9004.n50 a_2479_9004.n41 30.3012
R5728 a_2479_9004.n0 a_2479_9004.t3 28.5655
R5729 a_2479_9004.n0 a_2479_9004.t1 28.5655
R5730 a_2479_9004.t7 a_2479_9004.n72 28.5655
R5731 a_2479_9004.n72 a_2479_9004.t5 28.5655
R5732 a_2479_9004.n33 a_2479_9004.n9 24.8476
R5733 a_2479_9004.n64 a_2479_9004.n40 24.8476
R5734 a_2479_9004.n32 a_2479_9004.n16 23.3417
R5735 a_2479_9004.n63 a_2479_9004.n47 23.3417
R5736 a_2479_9004.n36 a_2479_9004.n35 22.0256
R5737 a_2479_9004.n67 a_2479_9004.n66 22.0256
R5738 a_2479_9004.n29 a_2479_9004.n15 21.8358
R5739 a_2479_9004.n60 a_2479_9004.n46 21.8358
R5740 a_2479_9004.n27 a_2479_9004.n14 20.3299
R5741 a_2479_9004.n58 a_2479_9004.n45 20.3299
R5742 a_2479_9004.n25 a_2479_9004.n13 18.824
R5743 a_2479_9004.n56 a_2479_9004.n44 18.824
R5744 a_2479_9004.n7 a_2479_9004.n5 17.4823
R5745 a_2479_9004.n23 a_2479_9004.n12 17.3181
R5746 a_2479_9004.n54 a_2479_9004.n43 17.3181
R5747 a_2479_9004.n34 a_2479_9004.n10 16.3559
R5748 a_2479_9004.n65 a_2479_9004.n41 16.3559
R5749 a_2479_9004.n21 a_2479_9004.n11 15.8123
R5750 a_2479_9004.n52 a_2479_9004.n42 15.8123
R5751 a_2479_9004.n7 a_2479_9004.n6 14.6053
R5752 a_2479_9004.n38 a_2479_9004.n37 14.377
R5753 a_2479_9004.n35 a_2479_9004.n9 12.7256
R5754 a_2479_9004.n66 a_2479_9004.n40 12.7256
R5755 a_2479_9004.n19 a_2479_9004.n11 11.2946
R5756 a_2479_9004.n50 a_2479_9004.n42 11.2946
R5757 a_2479_9004.n69 a_2479_9004.n7 10.4849
R5758 a_2479_9004.n21 a_2479_9004.n12 9.78874
R5759 a_2479_9004.n52 a_2479_9004.n43 9.78874
R5760 a_2479_9004.n9 a_2479_9004.n8 9.3005
R5761 a_2479_9004.n32 a_2479_9004.n31 9.3005
R5762 a_2479_9004.n30 a_2479_9004.n29 9.3005
R5763 a_2479_9004.n28 a_2479_9004.n27 9.3005
R5764 a_2479_9004.n26 a_2479_9004.n25 9.3005
R5765 a_2479_9004.n24 a_2479_9004.n23 9.3005
R5766 a_2479_9004.n22 a_2479_9004.n21 9.3005
R5767 a_2479_9004.n20 a_2479_9004.n19 9.3005
R5768 a_2479_9004.n40 a_2479_9004.n39 9.3005
R5769 a_2479_9004.n63 a_2479_9004.n62 9.3005
R5770 a_2479_9004.n61 a_2479_9004.n60 9.3005
R5771 a_2479_9004.n59 a_2479_9004.n58 9.3005
R5772 a_2479_9004.n57 a_2479_9004.n56 9.3005
R5773 a_2479_9004.n55 a_2479_9004.n54 9.3005
R5774 a_2479_9004.n53 a_2479_9004.n52 9.3005
R5775 a_2479_9004.n51 a_2479_9004.n50 9.3005
R5776 a_2479_9004.n70 a_2479_9004.n69 8.69704
R5777 a_2479_9004.n23 a_2479_9004.n13 8.28285
R5778 a_2479_9004.n54 a_2479_9004.n44 8.28285
R5779 a_2479_9004.n25 a_2479_9004.n14 6.77697
R5780 a_2479_9004.n56 a_2479_9004.n45 6.77697
R5781 a_2479_9004.n38 a_2479_9004.n36 6.19091
R5782 a_2479_9004.n27 a_2479_9004.n15 5.27109
R5783 a_2479_9004.n58 a_2479_9004.n46 5.27109
R5784 a_2479_9004.n29 a_2479_9004.n16 3.76521
R5785 a_2479_9004.n60 a_2479_9004.n47 3.76521
R5786 a_2479_9004.n68 a_2479_9004.n67 3.31388
R5787 a_2479_9004.n5 a_2479_9004.t16 2.48621
R5788 a_2479_9004.n5 a_2479_9004.t15 2.48621
R5789 a_2479_9004.n6 a_2479_9004.t20 2.48621
R5790 a_2479_9004.n6 a_2479_9004.t19 2.48621
R5791 a_2479_9004.n34 a_2479_9004.t17 2.48621
R5792 a_2479_9004.n34 a_2479_9004.t9 2.48621
R5793 a_2479_9004.n37 a_2479_9004.t14 2.48621
R5794 a_2479_9004.n37 a_2479_9004.t13 2.48621
R5795 a_2479_9004.n65 a_2479_9004.t12 2.48621
R5796 a_2479_9004.n65 a_2479_9004.t18 2.48621
R5797 a_2479_9004.n18 a_2479_9004.n10 2.36936
R5798 a_2479_9004.n49 a_2479_9004.n41 2.36936
R5799 a_2479_9004.n68 a_2479_9004.n38 2.30287
R5800 a_2479_9004.n33 a_2479_9004.n32 2.25932
R5801 a_2479_9004.n64 a_2479_9004.n63 2.25932
R5802 a_2479_9004.n69 a_2479_9004.n68 1.07418
R5803 a_2479_9004.n18 a_2479_9004.n17 0.320353
R5804 a_2479_9004.n49 a_2479_9004.n48 0.320353
R5805 a_2479_9004.n36 a_2479_9004.n8 0.196152
R5806 a_2479_9004.n31 a_2479_9004.n8 0.196152
R5807 a_2479_9004.n31 a_2479_9004.n30 0.196152
R5808 a_2479_9004.n30 a_2479_9004.n28 0.196152
R5809 a_2479_9004.n28 a_2479_9004.n26 0.196152
R5810 a_2479_9004.n26 a_2479_9004.n24 0.196152
R5811 a_2479_9004.n24 a_2479_9004.n22 0.196152
R5812 a_2479_9004.n22 a_2479_9004.n20 0.196152
R5813 a_2479_9004.n20 a_2479_9004.n18 0.196152
R5814 a_2479_9004.n67 a_2479_9004.n39 0.196152
R5815 a_2479_9004.n62 a_2479_9004.n39 0.196152
R5816 a_2479_9004.n62 a_2479_9004.n61 0.196152
R5817 a_2479_9004.n61 a_2479_9004.n59 0.196152
R5818 a_2479_9004.n59 a_2479_9004.n57 0.196152
R5819 a_2479_9004.n57 a_2479_9004.n55 0.196152
R5820 a_2479_9004.n55 a_2479_9004.n53 0.196152
R5821 a_2479_9004.n53 a_2479_9004.n51 0.196152
R5822 a_2479_9004.n51 a_2479_9004.n49 0.196152
R5823 a_2479_9004.n4 a_2479_9004.n3 0.0850588
R5824 a_2479_9004.n2 a_2479_9004.n1 0.0427794
R5825 a_2479_9004.n3 a_2479_9004.n2 0.0427794
R5826 a_2479_9004.n71 a_2479_9004.n4 0.0427794
R5827 a_2479_9004.n71 a_2479_9004.n70 0.0427794
R5828 a_3758_2896.n33 a_3758_2896.n32 185
R5829 a_3758_2896.n33 a_3758_2896.n15 185
R5830 a_3758_2896.n33 a_3758_2896.n14 185
R5831 a_3758_2896.n33 a_3758_2896.n13 185
R5832 a_3758_2896.n33 a_3758_2896.n12 185
R5833 a_3758_2896.n33 a_3758_2896.n11 185
R5834 a_3758_2896.n33 a_3758_2896.n10 185
R5835 a_3758_2896.n16 a_3758_2896.t13 130.75
R5836 a_3758_2896.n16 a_3758_2896.t14 91.3557
R5837 a_3758_2896.n34 a_3758_2896.n33 86.5152
R5838 a_3758_2896.n18 a_3758_2896.n9 30.3012
R5839 a_3758_2896.n2 a_3758_2896.n0 29.1073
R5840 a_3758_2896.n39 a_3758_2896.n38 27.9576
R5841 a_3758_2896.n37 a_3758_2896.n36 27.9576
R5842 a_3758_2896.n6 a_3758_2896.n5 27.9576
R5843 a_3758_2896.n4 a_3758_2896.n3 27.9576
R5844 a_3758_2896.n2 a_3758_2896.n1 27.9576
R5845 a_3758_2896.n32 a_3758_2896.n8 24.8476
R5846 a_3758_2896.n31 a_3758_2896.n15 23.3417
R5847 a_3758_2896.n35 a_3758_2896.n34 22.0256
R5848 a_3758_2896.n28 a_3758_2896.n14 21.8358
R5849 a_3758_2896.n26 a_3758_2896.n13 20.3299
R5850 a_3758_2896.n24 a_3758_2896.n12 18.824
R5851 a_3758_2896.n22 a_3758_2896.n11 17.3181
R5852 a_3758_2896.n33 a_3758_2896.n9 16.3559
R5853 a_3758_2896.n20 a_3758_2896.n10 15.8123
R5854 a_3758_2896.n34 a_3758_2896.n8 12.7256
R5855 a_3758_2896.n37 a_3758_2896.n35 12.0517
R5856 a_3758_2896.n18 a_3758_2896.n10 11.2946
R5857 a_3758_2896.n20 a_3758_2896.n11 9.78874
R5858 a_3758_2896.n8 a_3758_2896.n7 9.3005
R5859 a_3758_2896.n31 a_3758_2896.n30 9.3005
R5860 a_3758_2896.n29 a_3758_2896.n28 9.3005
R5861 a_3758_2896.n27 a_3758_2896.n26 9.3005
R5862 a_3758_2896.n25 a_3758_2896.n24 9.3005
R5863 a_3758_2896.n23 a_3758_2896.n22 9.3005
R5864 a_3758_2896.n21 a_3758_2896.n20 9.3005
R5865 a_3758_2896.n19 a_3758_2896.n18 9.3005
R5866 a_3758_2896.n22 a_3758_2896.n12 8.28285
R5867 a_3758_2896.n24 a_3758_2896.n13 6.77697
R5868 a_3758_2896.n36 a_3758_2896.t5 5.8005
R5869 a_3758_2896.n36 a_3758_2896.t7 5.8005
R5870 a_3758_2896.n5 a_3758_2896.t2 5.8005
R5871 a_3758_2896.n5 a_3758_2896.t1 5.8005
R5872 a_3758_2896.n3 a_3758_2896.t9 5.8005
R5873 a_3758_2896.n3 a_3758_2896.t8 5.8005
R5874 a_3758_2896.n1 a_3758_2896.t0 5.8005
R5875 a_3758_2896.n1 a_3758_2896.t10 5.8005
R5876 a_3758_2896.n0 a_3758_2896.t3 5.8005
R5877 a_3758_2896.n0 a_3758_2896.t4 5.8005
R5878 a_3758_2896.n39 a_3758_2896.t6 5.8005
R5879 a_3758_2896.t11 a_3758_2896.n39 5.8005
R5880 a_3758_2896.n26 a_3758_2896.n14 5.27109
R5881 a_3758_2896.n28 a_3758_2896.n15 3.76521
R5882 a_3758_2896.n33 a_3758_2896.t14 2.48621
R5883 a_3758_2896.n33 a_3758_2896.t12 2.48621
R5884 a_3758_2896.n17 a_3758_2896.n9 2.36936
R5885 a_3758_2896.n6 a_3758_2896.n4 2.30199
R5886 a_3758_2896.n32 a_3758_2896.n31 2.25932
R5887 a_3758_2896.n4 a_3758_2896.n2 1.1502
R5888 a_3758_2896.n38 a_3758_2896.n6 1.1502
R5889 a_3758_2896.n38 a_3758_2896.n37 1.1502
R5890 a_3758_2896.n17 a_3758_2896.n16 0.320353
R5891 a_3758_2896.n35 a_3758_2896.n7 0.196152
R5892 a_3758_2896.n30 a_3758_2896.n7 0.196152
R5893 a_3758_2896.n30 a_3758_2896.n29 0.196152
R5894 a_3758_2896.n29 a_3758_2896.n27 0.196152
R5895 a_3758_2896.n27 a_3758_2896.n25 0.196152
R5896 a_3758_2896.n25 a_3758_2896.n23 0.196152
R5897 a_3758_2896.n23 a_3758_2896.n21 0.196152
R5898 a_3758_2896.n21 a_3758_2896.n19 0.196152
R5899 a_3758_2896.n19 a_3758_2896.n17 0.196152
R5900 EN.n0 EN.t0 262.997
R5901 EN.n1 EN.t1 262.007
R5902 EN.n0 EN.t2 262.007
R5903 EN.n1 EN.n0 0.989232
R5904 EN EN.n1 0.365614
R5905 C1 C1.t0 17.7852
R5906 C1 C1.t1 0.00167066
R5907 IBIAS.n26 IBIAS.n25 185
R5908 IBIAS.n26 IBIAS.n8 185
R5909 IBIAS.n26 IBIAS.n7 185
R5910 IBIAS.n26 IBIAS.n6 185
R5911 IBIAS.n26 IBIAS.n5 185
R5912 IBIAS.n26 IBIAS.n4 185
R5913 IBIAS.n26 IBIAS.n3 185
R5914 IBIAS.n9 IBIAS.t0 130.75
R5915 IBIAS.n9 IBIAS.t1 91.3557
R5916 IBIAS.n27 IBIAS.n26 86.5152
R5917 IBIAS.n11 IBIAS.n2 30.3012
R5918 IBIAS.n25 IBIAS.n1 24.8476
R5919 IBIAS.n24 IBIAS.n8 23.3417
R5920 IBIAS.n28 IBIAS.n27 22.0256
R5921 IBIAS.n21 IBIAS.n7 21.8358
R5922 IBIAS.n19 IBIAS.n6 20.3299
R5923 IBIAS.n17 IBIAS.n5 18.824
R5924 IBIAS.n15 IBIAS.n4 17.3181
R5925 IBIAS.n26 IBIAS.n2 16.3559
R5926 IBIAS.n13 IBIAS.n3 15.8123
R5927 IBIAS.n27 IBIAS.n1 12.7256
R5928 IBIAS.n11 IBIAS.n3 11.2946
R5929 IBIAS.n13 IBIAS.n4 9.78874
R5930 IBIAS.n1 IBIAS.n0 9.3005
R5931 IBIAS.n24 IBIAS.n23 9.3005
R5932 IBIAS.n22 IBIAS.n21 9.3005
R5933 IBIAS.n20 IBIAS.n19 9.3005
R5934 IBIAS.n18 IBIAS.n17 9.3005
R5935 IBIAS.n16 IBIAS.n15 9.3005
R5936 IBIAS.n14 IBIAS.n13 9.3005
R5937 IBIAS.n12 IBIAS.n11 9.3005
R5938 IBIAS.n15 IBIAS.n5 8.28285
R5939 IBIAS.n17 IBIAS.n6 6.77697
R5940 IBIAS.n19 IBIAS.n7 5.27109
R5941 IBIAS IBIAS.n28 5.23142
R5942 IBIAS.n21 IBIAS.n8 3.76521
R5943 IBIAS.n26 IBIAS.t1 2.48621
R5944 IBIAS.n26 IBIAS.t2 2.48621
R5945 IBIAS.n10 IBIAS.n2 2.36936
R5946 IBIAS.n25 IBIAS.n24 2.25932
R5947 IBIAS.n10 IBIAS.n9 0.320353
R5948 IBIAS.n28 IBIAS.n0 0.196152
R5949 IBIAS.n23 IBIAS.n0 0.196152
R5950 IBIAS.n23 IBIAS.n22 0.196152
R5951 IBIAS.n22 IBIAS.n20 0.196152
R5952 IBIAS.n20 IBIAS.n18 0.196152
R5953 IBIAS.n18 IBIAS.n16 0.196152
R5954 IBIAS.n16 IBIAS.n14 0.196152
R5955 IBIAS.n14 IBIAS.n12 0.196152
R5956 IBIAS.n12 IBIAS.n10 0.196152
C0 VOUT VDD 9.72735f
C1 VOUT VN 0.15325f
C2 C1 VDD 0.11857f
C3 VOUT VP 0.4883f
C4 VN VP 5.95617f
C5 VOUT EN 0.69581f
C6 VOUT C1 57.8052f
C7 EN IBIAS 0.80152f
C8 IBIAS VSS 2.04035f
C9 EN VSS 3.05889f
C10 VP VSS 5.14937f
C11 VN VSS 5.45055f
C12 VOUT VSS 20.4866f
C13 VDD VSS 14.74629f
C14 C1 VSS 33.83365f
C15 C1.t0 VSS 0.2943f
C16 C1.t1 VSS 28.5579f
C17 a_3758_2896.t6 VSS 0.03416f
C18 a_3758_2896.t3 VSS 0.03416f
C19 a_3758_2896.t4 VSS 0.03416f
C20 a_3758_2896.n0 VSS 0.11734f
C21 a_3758_2896.t0 VSS 0.03416f
C22 a_3758_2896.t10 VSS 0.03416f
C23 a_3758_2896.n1 VSS 0.10037f
C24 a_3758_2896.n2 VSS 0.75156f
C25 a_3758_2896.t9 VSS 0.03416f
C26 a_3758_2896.t8 VSS 0.03416f
C27 a_3758_2896.n3 VSS 0.10037f
C28 a_3758_2896.n4 VSS 0.39548f
C29 a_3758_2896.t2 VSS 0.03416f
C30 a_3758_2896.t1 VSS 0.03416f
C31 a_3758_2896.n5 VSS 0.10037f
C32 a_3758_2896.n6 VSS 0.39548f
C33 a_3758_2896.n7 VSS 0.01301f
C34 a_3758_2896.t14 VSS 0.12182f
C35 a_3758_2896.n9 VSS 0.01076f
C36 a_3758_2896.t13 VSS 0.79281f
C37 a_3758_2896.n16 VSS 1.50323f
C38 a_3758_2896.n17 VSS 0.21382f
C39 a_3758_2896.n19 VSS 0.01301f
C40 a_3758_2896.n21 VSS 0.01301f
C41 a_3758_2896.n23 VSS 0.01301f
C42 a_3758_2896.n25 VSS 0.01301f
C43 a_3758_2896.n27 VSS 0.01301f
C44 a_3758_2896.n29 VSS 0.01301f
C45 a_3758_2896.n30 VSS 0.01301f
C46 a_3758_2896.t12 VSS 0.07972f
C47 a_3758_2896.n33 VSS 0.17055f
C48 a_3758_2896.n35 VSS 0.36219f
C49 a_3758_2896.t5 VSS 0.03416f
C50 a_3758_2896.t7 VSS 0.03416f
C51 a_3758_2896.n36 VSS 0.10037f
C52 a_3758_2896.n37 VSS 0.64652f
C53 a_3758_2896.n38 VSS 0.33874f
C54 a_3758_2896.n39 VSS 0.10037f
C55 a_3758_2896.t11 VSS 0.03416f
C56 a_2479_9004.t3 VSS 0.02166f
C57 a_2479_9004.t1 VSS 0.02166f
C58 a_2479_9004.n0 VSS 0.04534f
C59 a_2479_9004.t23 VSS 0.09411f
C60 a_2479_9004.t2 VSS 0.09411f
C61 a_2479_9004.n1 VSS -0.15502f
C62 a_2479_9004.n2 VSS 0.2387f
C63 a_2479_9004.t24 VSS 0.09411f
C64 a_2479_9004.t0 VSS 0.09411f
C65 a_2479_9004.n3 VSS 0.24905f
C66 a_2479_9004.t6 VSS 0.09411f
C67 a_2479_9004.t21 VSS 0.09411f
C68 a_2479_9004.n4 VSS 0.24905f
C69 a_2479_9004.t4 VSS 0.09411f
C70 a_2479_9004.t16 VSS 0.1516f
C71 a_2479_9004.t15 VSS 0.1516f
C72 a_2479_9004.n5 VSS 0.84136f
C73 a_2479_9004.t20 VSS 0.1516f
C74 a_2479_9004.t19 VSS 0.1516f
C75 a_2479_9004.n6 VSS 0.62542f
C76 a_2479_9004.n7 VSS 3.09987f
C77 a_2479_9004.n8 VSS 0.02473f
C78 a_2479_9004.n9 VSS 0.01699f
C79 a_2479_9004.t17 VSS 0.1516f
C80 a_2479_9004.n10 VSS 0.02047f
C81 a_2479_9004.t10 VSS 0.08006f
C82 a_2479_9004.t8 VSS 1.50795f
C83 a_2479_9004.n17 VSS 2.88661f
C84 a_2479_9004.n18 VSS 0.40663f
C85 a_2479_9004.n19 VSS 0.01649f
C86 a_2479_9004.n20 VSS 0.02473f
C87 a_2479_9004.n22 VSS 0.02473f
C88 a_2479_9004.n24 VSS 0.02473f
C89 a_2479_9004.n26 VSS 0.02473f
C90 a_2479_9004.n28 VSS 0.02473f
C91 a_2479_9004.n30 VSS 0.02473f
C92 a_2479_9004.n31 VSS 0.02473f
C93 a_2479_9004.t9 VSS 0.1516f
C94 a_2479_9004.n34 VSS 0.32433f
C95 a_2479_9004.n35 VSS 0.01069f
C96 a_2479_9004.n36 VSS 0.38075f
C97 a_2479_9004.t14 VSS 0.1516f
C98 a_2479_9004.t13 VSS 0.1516f
C99 a_2479_9004.n37 VSS 0.61041f
C100 a_2479_9004.n38 VSS 1.4281f
C101 a_2479_9004.n39 VSS 0.02473f
C102 a_2479_9004.n40 VSS 0.01699f
C103 a_2479_9004.t12 VSS 0.23166f
C104 a_2479_9004.n41 VSS 0.02047f
C105 a_2479_9004.t11 VSS 1.50795f
C106 a_2479_9004.n48 VSS 2.88661f
C107 a_2479_9004.n49 VSS 0.40663f
C108 a_2479_9004.n50 VSS 0.01649f
C109 a_2479_9004.n51 VSS 0.02473f
C110 a_2479_9004.n53 VSS 0.02473f
C111 a_2479_9004.n55 VSS 0.02473f
C112 a_2479_9004.n57 VSS 0.02473f
C113 a_2479_9004.n59 VSS 0.02473f
C114 a_2479_9004.n61 VSS 0.02473f
C115 a_2479_9004.n62 VSS 0.02473f
C116 a_2479_9004.t18 VSS 0.1516f
C117 a_2479_9004.n65 VSS 0.32433f
C118 a_2479_9004.n66 VSS 0.01069f
C119 a_2479_9004.n67 VSS 0.19498f
C120 a_2479_9004.n68 VSS 0.36196f
C121 a_2479_9004.n69 VSS 1.87446f
C122 a_2479_9004.t22 VSS 0.09411f
C123 a_2479_9004.n70 VSS 0.94824f
C124 a_2479_9004.n71 VSS 0.2387f
C125 a_2479_9004.t5 VSS 0.02166f
C126 a_2479_9004.n72 VSS 0.04534f
C127 a_2479_9004.t7 VSS 0.02166f
C128 VN.t0 VSS 1.38469f
C129 VN.t1 VSS 1.38075f
C130 VN.n0 VSS 1.21869f
C131 VN.t4 VSS 1.38075f
C132 VN.n1 VSS 0.60854f
C133 VN.t5 VSS 1.38202f
C134 VN.n2 VSS 1.32742f
C135 VN.t7 VSS 1.38043f
C136 VN.t2 VSS 1.38365f
C137 VN.t6 VSS 1.38043f
C138 VN.n3 VSS 1.20405f
C139 VN.n4 VSS 0.57632f
C140 VN.t3 VSS 1.38021f
C141 VN.n5 VSS 0.59805f
C142 VN.n6 VSS 0.73649f
C143 a_2995_7336.t10 VSS 0.11279f
C144 a_2995_7336.t1 VSS 0.11279f
C145 a_2995_7336.n0 VSS 0.32268f
C146 a_2995_7336.t18 VSS 0.11279f
C147 a_2995_7336.t11 VSS 0.11279f
C148 a_2995_7336.n1 VSS 0.32268f
C149 a_2995_7336.t12 VSS 0.11279f
C150 a_2995_7336.t4 VSS 0.11279f
C151 a_2995_7336.n2 VSS 0.32272f
C152 a_2995_7336.n3 VSS 1.26812f
C153 a_2995_7336.n4 VSS 0.0184f
C154 a_2995_7336.n5 VSS 0.01264f
C155 a_2995_7336.t2 VSS 0.11279f
C156 a_2995_7336.n6 VSS 0.01523f
C157 a_2995_7336.t7 VSS 0.05957f
C158 a_2995_7336.t5 VSS 1.12173f
C159 a_2995_7336.n13 VSS 2.1269f
C160 a_2995_7336.n14 VSS 0.30254f
C161 a_2995_7336.n15 VSS 0.01227f
C162 a_2995_7336.n16 VSS 0.0184f
C163 a_2995_7336.n18 VSS 0.0184f
C164 a_2995_7336.n20 VSS 0.0184f
C165 a_2995_7336.n22 VSS 0.0184f
C166 a_2995_7336.n24 VSS 0.0184f
C167 a_2995_7336.n26 VSS 0.0184f
C168 a_2995_7336.n27 VSS 0.0184f
C169 a_2995_7336.t6 VSS 0.11279f
C170 a_2995_7336.n30 VSS 0.24131f
C171 a_2995_7336.n32 VSS 0.18922f
C172 a_2995_7336.t19 VSS 0.11279f
C173 a_2995_7336.t16 VSS 0.11279f
C174 a_2995_7336.n33 VSS 0.32268f
C175 a_2995_7336.t17 VSS 0.11279f
C176 a_2995_7336.t9 VSS 0.11279f
C177 a_2995_7336.n34 VSS 0.32272f
C178 a_2995_7336.t15 VSS 0.11279f
C179 a_2995_7336.t3 VSS 0.11279f
C180 a_2995_7336.n35 VSS 0.32268f
C181 a_2995_7336.t8 VSS 0.11279f
C182 a_2995_7336.t13 VSS 0.11279f
C183 a_2995_7336.n36 VSS 0.32272f
C184 a_2995_7336.n37 VSS 1.26812f
C185 a_2995_7336.n38 VSS 1.58502f
C186 a_2995_7336.n39 VSS 1.93909f
C187 a_2995_7336.n40 VSS 1.60511f
C188 a_2995_7336.t14 VSS 0.11279f
C189 a_2995_7336.n41 VSS 0.32269f
C190 a_2995_7336.t0 VSS 0.11279f
C191 VP.t7 VSS 1.38738f
C192 VP.t6 VSS 1.38343f
C193 VP.n0 VSS 1.22106f
C194 VP.t2 VSS 1.38343f
C195 VP.n1 VSS 0.60972f
C196 VP.t1 VSS 1.3847f
C197 VP.n2 VSS 1.27437f
C198 VP.t3 VSS 1.38633f
C199 VP.t5 VSS 1.38311f
C200 VP.n3 VSS 1.20639f
C201 VP.t4 VSS 1.38311f
C202 VP.n4 VSS 0.57744f
C203 VP.t0 VSS 1.38289f
C204 VP.n5 VSS 0.59921f
C205 VP.n6 VSS 0.717f
C206 a_4920_2896.t10 VSS 0.02015f
C207 a_4920_2896.t16 VSS 0.02015f
C208 a_4920_2896.n0 VSS 0.04651f
C209 a_4920_2896.t4 VSS 0.02015f
C210 a_4920_2896.t11 VSS 0.02015f
C211 a_4920_2896.n1 VSS 0.04651f
C212 a_4920_2896.t20 VSS 0.02015f
C213 a_4920_2896.t3 VSS 0.02015f
C214 a_4920_2896.n2 VSS 0.04651f
C215 a_4920_2896.t22 VSS 0.02015f
C216 a_4920_2896.t21 VSS 0.02015f
C217 a_4920_2896.n3 VSS 0.04651f
C218 a_4920_2896.t14 VSS 0.02015f
C219 a_4920_2896.t9 VSS 0.02015f
C220 a_4920_2896.n4 VSS 0.05823f
C221 a_4920_2896.n5 VSS 0.44309f
C222 a_4920_2896.n6 VSS 0.18382f
C223 a_4920_2896.n7 VSS 0.18382f
C224 a_4920_2896.n8 VSS 0.18382f
C225 a_4920_2896.t8 VSS 0.02015f
C226 a_4920_2896.t1 VSS 0.02015f
C227 a_4920_2896.n9 VSS 0.04759f
C228 a_4920_2896.t18 VSS 0.02015f
C229 a_4920_2896.t2 VSS 0.02015f
C230 a_4920_2896.n10 VSS 0.04759f
C231 a_4920_2896.t13 VSS 0.02015f
C232 a_4920_2896.t19 VSS 0.02015f
C233 a_4920_2896.n11 VSS 0.04759f
C234 a_4920_2896.t5 VSS 0.02015f
C235 a_4920_2896.t12 VSS 0.02015f
C236 a_4920_2896.n12 VSS 0.04759f
C237 a_4920_2896.t7 VSS 0.02015f
C238 a_4920_2896.t6 VSS 0.02015f
C239 a_4920_2896.n13 VSS 0.04759f
C240 a_4920_2896.t0 VSS 0.02015f
C241 a_4920_2896.t17 VSS 0.02015f
C242 a_4920_2896.n14 VSS 0.05955f
C243 a_4920_2896.n15 VSS 0.4586f
C244 a_4920_2896.n16 VSS 0.1917f
C245 a_4920_2896.n17 VSS 0.1917f
C246 a_4920_2896.n18 VSS 0.1917f
C247 a_4920_2896.n19 VSS 0.37064f
C248 a_4920_2896.t26 VSS 0.07185f
C249 a_4920_2896.t25 VSS 0.46761f
C250 a_4920_2896.n30 VSS 0.88664f
C251 a_4920_2896.n44 VSS 0.12612f
C252 a_4920_2896.t24 VSS 0.04702f
C253 a_4920_2896.n46 VSS 0.10059f
C254 a_4920_2896.n48 VSS 0.0652f
C255 a_4920_2896.n49 VSS 0.31283f
C256 a_4920_2896.n50 VSS 0.23403f
C257 a_4920_2896.t15 VSS 0.02015f
C258 a_4920_2896.n51 VSS 0.04651f
C259 a_4920_2896.t23 VSS 0.02015f
C260 a_2080_2896.t7 VSS 0.02936f
C261 a_2080_2896.t22 VSS 0.21364f
C262 a_2080_2896.t30 VSS 0.21316f
C263 a_2080_2896.n9 VSS 0.22163f
C264 a_2080_2896.t9 VSS 0.21316f
C265 a_2080_2896.n10 VSS 0.08384f
C266 a_2080_2896.t10 VSS 0.21316f
C267 a_2080_2896.n11 VSS 0.08384f
C268 a_2080_2896.t11 VSS 0.21316f
C269 a_2080_2896.n12 VSS 0.08384f
C270 a_2080_2896.t40 VSS 0.21316f
C271 a_2080_2896.n13 VSS 0.08384f
C272 a_2080_2896.t39 VSS 0.21316f
C273 a_2080_2896.n14 VSS 0.08384f
C274 a_2080_2896.t28 VSS 0.21316f
C275 a_2080_2896.n15 VSS 0.08384f
C276 a_2080_2896.t29 VSS 0.21316f
C277 a_2080_2896.n16 VSS 0.08384f
C278 a_2080_2896.t18 VSS 0.21316f
C279 a_2080_2896.n17 VSS 0.08384f
C280 a_2080_2896.t8 VSS 0.21316f
C281 a_2080_2896.n18 VSS 0.08384f
C282 a_2080_2896.t21 VSS 0.21316f
C283 a_2080_2896.n19 VSS 0.11277f
C284 a_2080_2896.t35 VSS 0.21356f
C285 a_2080_2896.t43 VSS 0.21238f
C286 a_2080_2896.t27 VSS 0.21229f
C287 a_2080_2896.n20 VSS 0.1205f
C288 a_2080_2896.n21 VSS 0.13801f
C289 a_2080_2896.t15 VSS 0.21238f
C290 a_2080_2896.t38 VSS 0.21229f
C291 a_2080_2896.n22 VSS 0.1205f
C292 a_2080_2896.n23 VSS 0.02104f
C293 a_2080_2896.t32 VSS 0.21238f
C294 a_2080_2896.t16 VSS 0.21229f
C295 a_2080_2896.n24 VSS 0.1205f
C296 a_2080_2896.n25 VSS 0.02104f
C297 a_2080_2896.t33 VSS 0.21238f
C298 a_2080_2896.t17 VSS 0.21229f
C299 a_2080_2896.n26 VSS 0.1205f
C300 a_2080_2896.n27 VSS 0.02104f
C301 a_2080_2896.t34 VSS 0.21238f
C302 a_2080_2896.t19 VSS 0.21229f
C303 a_2080_2896.n28 VSS 0.1205f
C304 a_2080_2896.n29 VSS 0.02104f
C305 a_2080_2896.n30 VSS 0.02104f
C306 a_2080_2896.t23 VSS 0.21238f
C307 a_2080_2896.n31 VSS 0.01136f
C308 a_2080_2896.t25 VSS 0.21238f
C309 a_2080_2896.n32 VSS 0.07247f
C310 a_2080_2896.n33 VSS 0.04758f
C311 a_2080_2896.t5 VSS 0.16153f
C312 a_2080_2896.t6 VSS 0.01258f
C313 a_2080_2896.t4 VSS 0.01258f
C314 a_2080_2896.n53 VSS 0.02517f
C315 a_2080_2896.n56 VSS 0.11181f
C316 a_2080_2896.t3 VSS 0.16153f
C317 a_2080_2896.n57 VSS 0.04758f
C318 a_2080_2896.n58 VSS 0.07247f
C319 a_2080_2896.n59 VSS 0.02104f
C320 a_2080_2896.t12 VSS 0.21238f
C321 a_2080_2896.t36 VSS 0.21229f
C322 a_2080_2896.n60 VSS 0.1205f
C323 a_2080_2896.n61 VSS 0.02104f
C324 a_2080_2896.t13 VSS 0.21238f
C325 a_2080_2896.t37 VSS 0.21229f
C326 a_2080_2896.n62 VSS 0.1205f
C327 a_2080_2896.n63 VSS 0.02104f
C328 a_2080_2896.t41 VSS 0.21238f
C329 a_2080_2896.t24 VSS 0.21229f
C330 a_2080_2896.n64 VSS 0.1205f
C331 a_2080_2896.n65 VSS 0.02104f
C332 a_2080_2896.t31 VSS 0.21238f
C333 a_2080_2896.t14 VSS 0.21229f
C334 a_2080_2896.n66 VSS 0.1205f
C335 a_2080_2896.n67 VSS 0.02104f
C336 a_2080_2896.t42 VSS 0.21238f
C337 a_2080_2896.t26 VSS 0.21229f
C338 a_2080_2896.n68 VSS 0.1205f
C339 a_2080_2896.n69 VSS 0.02104f
C340 a_2080_2896.t20 VSS 0.21316f
C341 a_2080_2896.n70 VSS 0.16653f
C342 a_2080_2896.n71 VSS 0.2988f
C343 a_2080_2896.n72 VSS 0.17452f
C344 a_2080_2896.t1 VSS 0.02936f
C345 a_2080_2896.n86 VSS 0.06282f
C346 a_2080_2896.n90 VSS 0.07876f
C347 a_2080_2896.t0 VSS 0.29202f
C348 a_2080_2896.n91 VSS 0.47059f
C349 a_2080_2896.n92 VSS 0.08427f
C350 a_2080_2896.t2 VSS 0.01433f
C351 VDD.t23 VSS 0.03729f
C352 VDD.t68 VSS 0.01296f
C353 VDD.n0 VSS 0.01158f
C354 VDD.t21 VSS 0.03444f
C355 VDD.n1 VSS 0.20115f
C356 VDD.n2 VSS 0.01756f
C357 VDD.n3 VSS 0.18618f
C358 VDD.n4 VSS 0.01756f
C359 VDD.n5 VSS 0.12574f
C360 VDD.n6 VSS 0.01756f
C361 VDD.n7 VSS 0.12574f
C362 VDD.n8 VSS 0.01756f
C363 VDD.n9 VSS 0.16718f
C364 VDD.n10 VSS 0.05232f
C365 VDD.t17 VSS 0.01585f
C366 VDD.n11 VSS 0.02495f
C367 VDD.n12 VSS 0.02539f
C368 VDD.t29 VSS 0.03447f
C369 VDD.t40 VSS 0.06759f
C370 VDD.t41 VSS 0.03736f
C371 VDD.n13 VSS 0.04502f
C372 VDD.n14 VSS 0.01651f
C373 VDD.n15 VSS 0.0203f
C374 VDD.n16 VSS 0.07594f
C375 VDD.n17 VSS 0.04082f
C376 VDD.t15 VSS 0.06755f
C377 VDD.n18 VSS 0.02539f
C378 VDD.n19 VSS 0.04082f
C379 VDD.t51 VSS 0.06757f
C380 VDD.n20 VSS 0.05959f
C381 VDD.n21 VSS 0.01946f
C382 VDD.n22 VSS 0.0203f
C383 VDD.n23 VSS 0.01651f
C384 VDD.t53 VSS 0.01585f
C385 VDD.n24 VSS 0.01653f
C386 VDD.t31 VSS 0.01585f
C387 VDD.n25 VSS 0.01653f
C388 VDD.n26 VSS 0.10792f
C389 VDD.n27 VSS 0.01756f
C390 VDD.n28 VSS 0.24218f
C391 VDD.n29 VSS 0.05232f
C392 VDD.n30 VSS 0.0203f
C393 VDD.t14 VSS 0.02943f
C394 VDD.n31 VSS 0.07594f
C395 VDD.n32 VSS 0.02539f
C396 VDD.t54 VSS 0.03447f
C397 VDD.n33 VSS 0.01946f
C398 VDD.n34 VSS 0.05959f
C399 VDD.t32 VSS 0.06757f
C400 VDD.n35 VSS 0.02495f
C401 VDD.n36 VSS 0.04082f
C402 VDD.t35 VSS 0.06755f
C403 VDD.n37 VSS 0.02539f
C404 VDD.n38 VSS 0.04082f
C405 VDD.t11 VSS 0.06759f
C406 VDD.n39 VSS 0.04502f
C407 VDD.n40 VSS 0.0203f
C408 VDD.n41 VSS 0.01651f
C409 VDD.t37 VSS 0.01585f
C410 VDD.n42 VSS 0.01651f
C411 VDD.t34 VSS 0.01585f
C412 VDD.n43 VSS 0.01653f
C413 VDD.t55 VSS 0.01585f
C414 VDD.n44 VSS 0.01653f
C415 VDD.n45 VSS 0.08183f
C416 VDD.n46 VSS 0.07903f
C417 VDD.n47 VSS 0.0311f
C418 VDD.n48 VSS 0.09167f
C419 VDD.n53 VSS 0.52396f
C420 VDD.n64 VSS 0.01365f
C421 VDD.n67 VSS 0.01329f
C422 VDD.n70 VSS 0.36362f
C423 VDD.n72 VSS 0.01329f
C424 VDD.n75 VSS 0.36935f
C425 VDD.t36 VSS 0.1947f
C426 VDD.n79 VSS 0.37508f
C427 VDD.n83 VSS 0.3808f
C428 VDD.t19 VSS 0.1947f
C429 VDD.n87 VSS 0.38653f
C430 VDD.n91 VSS 0.38939f
C431 VDD.t4 VSS 0.1947f
C432 VDD.t2 VSS 0.1947f
C433 VDD.t0 VSS 0.1947f
C434 VDD.n98 VSS 0.38653f
C435 VDD.t30 VSS 0.1947f
C436 VDD.t52 VSS 0.1947f
C437 VDD.n105 VSS 0.37508f
C438 VDD.t16 VSS 0.1947f
C439 VDD.n110 VSS 0.01329f
C440 VDD.n111 VSS 0.01329f
C441 VDD.t22 VSS 0.1947f
C442 VDD.n112 VSS 0.36362f
C443 VDD.n113 VSS 0.01329f
C444 VDD.n115 VSS 0.52396f
C445 VDD.n116 VSS 0.66426f
C446 VDD.n139 VSS 0.01365f
C447 VDD.n140 VSS 0.01365f
C448 VDD.n149 VSS 0.09305f
C449 VDD.n172 VSS 0.09305f
C450 VDD.n187 VSS 0.01365f
C451 VDD.n188 VSS 0.01365f
C452 VDD.n189 VSS 0.01329f
C453 VDD.n192 VSS 0.22619f
C454 VDD.n198 VSS 0.36935f
C455 VDD.n199 VSS 0.22046f
C456 VDD.n205 VSS 0.21474f
C457 VDD.n211 VSS 0.3808f
C458 VDD.n212 VSS 0.20901f
C459 VDD.n218 VSS 0.20329f
C460 VDD.n224 VSS 0.19756f
C461 VDD.n230 VSS 0.19756f
C462 VDD.t8 VSS 0.1947f
C463 VDD.n236 VSS 0.20329f
C464 VDD.n242 VSS 0.20901f
C465 VDD.t33 VSS 0.1947f
C466 VDD.n248 VSS 0.21474f
C467 VDD.n254 VSS 0.22046f
C468 VDD.n290 VSS 0.01365f
C469 VDD.n291 VSS 0.01329f
C470 VDD.t12 VSS 0.1947f
C471 VDD.n294 VSS 0.22619f
C472 VDD.n297 VSS 0.01329f
C473 VDD.n308 VSS 0.09401f
C474 VDD.n311 VSS 0.01365f
C475 VDD.n312 VSS 0.01365f
C476 VDD.n314 VSS 0.66426f
C477 VDD.n319 VSS 0.03228f
C478 VDD.n320 VSS 0.02337f
C479 VDD.n321 VSS 0.07085f
C480 VDD.n322 VSS 0.05232f
C481 VDD.t28 VSS 0.01585f
C482 VDD.n323 VSS 0.01946f
C483 VDD.n324 VSS 0.07594f
C484 VDD.n325 VSS 0.04082f
C485 VDD.t49 VSS 0.06759f
C486 VDD.t50 VSS 0.03736f
C487 VDD.n326 VSS 0.01651f
C488 VDD.n327 VSS 0.0203f
C489 VDD.n328 VSS 0.04502f
C490 VDD.n329 VSS 0.02539f
C491 VDD.t27 VSS 0.06755f
C492 VDD.n330 VSS 0.02539f
C493 VDD.t38 VSS 0.03447f
C494 VDD.n331 VSS 0.05959f
C495 VDD.t56 VSS 0.06757f
C496 VDD.n332 VSS 0.04082f
C497 VDD.n333 VSS 0.02495f
C498 VDD.n334 VSS 0.0203f
C499 VDD.n335 VSS 0.01651f
C500 VDD.t57 VSS 0.01585f
C501 VDD.n336 VSS 0.01653f
C502 VDD.t39 VSS 0.01585f
C503 VDD.n337 VSS 0.01653f
C504 VDD.n338 VSS 0.10809f
C505 VDD.n339 VSS 0.01756f
C506 VDD.n340 VSS 0.24293f
C507 VDD.n341 VSS 0.05232f
C508 VDD.n342 VSS 0.0203f
C509 VDD.n343 VSS 0.04502f
C510 VDD.n344 VSS 0.02495f
C511 VDD.t26 VSS 0.02943f
C512 VDD.n345 VSS 0.04082f
C513 VDD.t18 VSS 0.03447f
C514 VDD.t42 VSS 0.06757f
C515 VDD.n346 VSS 0.05959f
C516 VDD.n347 VSS 0.01946f
C517 VDD.n348 VSS 0.02539f
C518 VDD.t47 VSS 0.06755f
C519 VDD.n349 VSS 0.02539f
C520 VDD.t24 VSS 0.06759f
C521 VDD.n350 VSS 0.04082f
C522 VDD.n351 VSS 0.07594f
C523 VDD.n352 VSS 0.0203f
C524 VDD.n353 VSS 0.01651f
C525 VDD.t48 VSS 0.01585f
C526 VDD.n354 VSS 0.01651f
C527 VDD.t43 VSS 0.01585f
C528 VDD.n355 VSS 0.01653f
C529 VDD.t20 VSS 0.01585f
C530 VDD.n356 VSS 0.01653f
C531 VDD.n357 VSS 0.08183f
C532 VDD.n358 VSS 0.09923f
C533 VDD.n359 VSS 0.01814f
C534 VDD.n360 VSS 0.01756f
C535 VDD.n361 VSS 0.32081f
C536 VDD.n362 VSS 0.01756f
C537 VDD.n363 VSS 0.12574f
C538 VDD.n364 VSS 0.01756f
C539 VDD.n365 VSS 0.12574f
C540 VDD.t46 VSS 0.02937f
C541 VDD.n366 VSS 0.01653f
C542 VDD.n367 VSS 0.11223f
C543 VDD.t44 VSS 0.03444f
C544 VDD.n368 VSS 0.07391f
C545 VDD.n369 VSS 0.10272f
C546 VDD.n370 VSS 0.41333f
C547 VDD.n371 VSS 0.26414f
C548 VDD.n372 VSS 0.19973f
C549 VOUT.n0 VSS 0.01561f
C550 VOUT.n1 VSS 0.01513f
C551 VOUT.n2 VSS 0.2765f
C552 VOUT.n3 VSS 0.01513f
C553 VOUT.n4 VSS 0.11605f
C554 VOUT.n5 VSS 0.01513f
C555 VOUT.n6 VSS 0.11605f
C556 VOUT.n7 VSS 0.03194f
C557 VOUT.n8 VSS 0.03838f
C558 VOUT.t8 VSS 0.05763f
C559 VOUT.t10 VSS 0.02509f
C560 VOUT.n9 VSS 0.01408f
C561 VOUT.t5 VSS 0.01351f
C562 VOUT.n10 VSS 0.01408f
C563 VOUT.n11 VSS 0.01731f
C564 VOUT.n12 VSS 0.06898f
C565 VOUT.n13 VSS 0.0566f
C566 VOUT.t4 VSS 0.05761f
C567 VOUT.n14 VSS 0.02164f
C568 VOUT.n15 VSS 0.04613f
C569 VOUT.n16 VSS 0.10296f
C570 VOUT.t0 VSS 0.04729f
C571 VOUT.t13 VSS 0.02497f
C572 VOUT.t11 VSS 0.47028f
C573 VOUT.n26 VSS 0.89169f
C574 VOUT.n27 VSS 0.12684f
C575 VOUT.t12 VSS 0.04729f
C576 VOUT.n43 VSS 0.10117f
C577 VOUT.n45 VSS 0.44202f
C578 VOUT.n46 VSS 0.66145f
C579 VOUT.n48 VSS 0.01789f
C580 VOUT.t1 VSS 66.8769f
C581 VOUT.n49 VSS 0.03885f
C582 VOUT.n50 VSS 0.03489f
C583 VOUT.n51 VSS 1.16187f
C584 VOUT.n52 VSS 0.02957f
C585 VOUT.n53 VSS 0.02031f
C586 VOUT.n54 VSS 0.02041f
C587 VOUT.n55 VSS 0.06898f
C588 VOUT.t3 VSS 0.03185f
C589 VOUT.t6 VSS 0.05761f
C590 VOUT.n56 VSS 0.0566f
C591 VOUT.t2 VSS 0.05763f
C592 VOUT.n57 VSS 0.03838f
C593 VOUT.n58 VSS 0.01731f
C594 VOUT.n59 VSS 0.01408f
C595 VOUT.t7 VSS 0.01351f
C596 VOUT.n60 VSS 0.01408f
C597 VOUT.n61 VSS 0.0334f
C598 VOUT.n62 VSS 0.06133f
C599 VOUT.n63 VSS 0.01513f
C600 VOUT.n64 VSS 0.18517f
C601 VOUT.n65 VSS 0.01513f
C602 VOUT.n66 VSS 0.11605f
C603 VOUT.n67 VSS 0.01513f
C604 VOUT.n68 VSS 0.11605f
C605 VOUT.n69 VSS 0.01513f
C606 VOUT.n70 VSS 0.16056f
C607 VOUT.n71 VSS 0.27023f
C608 VOUT.n72 VSS 0.3823f
C609 a_2479_7336.t31 VSS 0.07294f
C610 a_2479_7336.t22 VSS 0.07285f
C611 a_2479_7336.n0 VSS 0.13526f
C612 a_2479_7336.t24 VSS 0.07285f
C613 a_2479_7336.n1 VSS 0.06289f
C614 a_2479_7336.n2 VSS 0.01915f
C615 a_2479_7336.n3 VSS 0.01315f
C616 a_2479_7336.t15 VSS 0.17933f
C617 a_2479_7336.n11 VSS 0.01276f
C618 a_2479_7336.t14 VSS 1.16729f
C619 a_2479_7336.n12 VSS 2.2345f
C620 a_2479_7336.n14 VSS 0.01915f
C621 a_2479_7336.n16 VSS 0.01915f
C622 a_2479_7336.n18 VSS 0.01915f
C623 a_2479_7336.n20 VSS 0.01915f
C624 a_2479_7336.n22 VSS 0.01915f
C625 a_2479_7336.n24 VSS 0.01915f
C626 a_2479_7336.n25 VSS 0.01915f
C627 a_2479_7336.n26 VSS 0.31477f
C628 a_2479_7336.n27 VSS 0.01585f
C629 a_2479_7336.t6 VSS 0.11735f
C630 a_2479_7336.n28 VSS 0.25106f
C631 a_2479_7336.n30 VSS 0.29467f
C632 a_2479_7336.t1 VSS 0.11735f
C633 a_2479_7336.t7 VSS 0.11735f
C634 a_2479_7336.n31 VSS 0.47249f
C635 a_2479_7336.n32 VSS 1.10557f
C636 a_2479_7336.n33 VSS 0.01915f
C637 a_2479_7336.n34 VSS 0.01315f
C638 a_2479_7336.t5 VSS 0.11735f
C639 a_2479_7336.n42 VSS 0.01276f
C640 a_2479_7336.t13 VSS 0.06198f
C641 a_2479_7336.t11 VSS 1.16729f
C642 a_2479_7336.n43 VSS 2.2345f
C643 a_2479_7336.n45 VSS 0.01915f
C644 a_2479_7336.n47 VSS 0.01915f
C645 a_2479_7336.n49 VSS 0.01915f
C646 a_2479_7336.n51 VSS 0.01915f
C647 a_2479_7336.n53 VSS 0.01915f
C648 a_2479_7336.n55 VSS 0.01915f
C649 a_2479_7336.n56 VSS 0.01915f
C650 a_2479_7336.n57 VSS 0.31477f
C651 a_2479_7336.n58 VSS 0.01585f
C652 a_2479_7336.t12 VSS 0.11735f
C653 a_2479_7336.n59 VSS 0.25106f
C654 a_2479_7336.n61 VSS 0.15093f
C655 a_2479_7336.n62 VSS 1.05081f
C656 a_2479_7336.t16 VSS 0.11735f
C657 a_2479_7336.t17 VSS 0.11735f
C658 a_2479_7336.n63 VSS 0.48416f
C659 a_2479_7336.n64 VSS 1.62989f
C660 a_2479_7336.t4 VSS 0.11735f
C661 a_2479_7336.t3 VSS 0.11735f
C662 a_2479_7336.n65 VSS 0.48416f
C663 a_2479_7336.n66 VSS 1.46324f
C664 a_2479_7336.t10 VSS 0.01676f
C665 a_2479_7336.t8 VSS 0.01676f
C666 a_2479_7336.n67 VSS 0.03536f
C667 a_2479_7336.t19 VSS 0.07294f
C668 a_2479_7336.t28 VSS 0.07285f
C669 a_2479_7336.n68 VSS 0.13526f
C670 a_2479_7336.t35 VSS 0.07285f
C671 a_2479_7336.n69 VSS 0.06289f
C672 a_2479_7336.n70 VSS 0.16351f
C673 a_2479_7336.t32 VSS 0.07285f
C674 a_2479_7336.n71 VSS 0.06289f
C675 a_2479_7336.t26 VSS 0.07285f
C676 a_2479_7336.n72 VSS 0.07206f
C677 a_2479_7336.t23 VSS 0.07285f
C678 a_2479_7336.n73 VSS 0.07206f
C679 a_2479_7336.t20 VSS 0.07285f
C680 a_2479_7336.n74 VSS 0.07206f
C681 a_2479_7336.t30 VSS 0.07285f
C682 a_2479_7336.n75 VSS 0.07206f
C683 a_2479_7336.t25 VSS 0.07285f
C684 a_2479_7336.n76 VSS 0.12272f
C685 a_2479_7336.t9 VSS 0.72083f
C686 a_2479_7336.n77 VSS 5.01204f
C687 a_2479_7336.n78 VSS 2.28905f
C688 a_2479_7336.t34 VSS 0.07285f
C689 a_2479_7336.n79 VSS 0.12615f
C690 a_2479_7336.t21 VSS 0.07285f
C691 a_2479_7336.n80 VSS 0.07206f
C692 a_2479_7336.t29 VSS 0.07285f
C693 a_2479_7336.n81 VSS 0.07206f
C694 a_2479_7336.t18 VSS 0.07285f
C695 a_2479_7336.n82 VSS 0.07206f
C696 a_2479_7336.t33 VSS 0.07285f
C697 a_2479_7336.n83 VSS 0.07206f
C698 a_2479_7336.t27 VSS 0.07285f
C699 a_2479_7336.n84 VSS 0.06289f
C700 a_2479_7336.n85 VSS 0.16351f
C701 a_2479_7336.t2 VSS 0.01676f
C702 a_2479_7336.n86 VSS 0.03536f
C703 a_2479_7336.t0 VSS 0.01676f
.ends

