* NGSPICE file created from ttsky25_two_stage_opamp.ext - technology: sky130A

.subckt ttsky25_two_stage_opamp VDD IBIAS VOUT VN VP EN VSS
X0 VSS.t132 VSS.t131 VSS.t132 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X1 VDD.t74 a_2479_7336.t18 VOUT.t26 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X2 VSS.t58 a_2080_2896.t5 a_2080_2896.t6 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X3 VDD.t73 a_2479_7336.t19 VOUT.t24 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X4 VDD.t55 VDD.t54 VDD.t55 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X5 VSS.t39 a_2080_2896.t8 a_4920_2896.t23 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 VSS.t17 a_2080_2896.t9 a_4920_2896.t22 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X7 a_2479_7336.t14 a_2479_7336.t13 a_2479_7336.t14 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X8 VSS.t130 VSS.t129 VSS.t130 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X9 VDD.t53 VDD.t52 VDD.t53 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X10 VDD.t72 a_2479_7336.t20 VOUT.t25 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X11 VDD.t71 a_2479_7336.t21 VOUT.t18 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X12 a_4920_2896.t21 a_2080_2896.t10 VSS.t64 VSS.t53 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X13 a_2479_7336.t12 a_2479_7336.t10 a_2479_7336.t11 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X14 a_2479_7336.t7 VP.t0 a_2995_7336.t14 VSS.t43 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X15 VSS.t56 a_2080_2896.t11 a_4920_2896.t20 VSS.t55 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 VSS.t128 VSS.t127 VSS.t128 VSS.t91 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X17 a_2995_7336.t2 VN.t0 a_2479_9004.t20 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X18 VDD.t70 a_2479_7336.t22 VOUT.t15 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X19 a_2479_9004.t19 VN.t1 a_2995_7336.t6 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X20 VSS.t126 VSS.t125 VSS.t126 VSS.t88 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X21 a_2479_9004.t12 a_2479_9004.t11 a_2479_9004.t12 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X22 VSS.t124 VSS.t123 VSS.t124 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X23 a_4920_2896.t19 a_2080_2896.t12 VSS.t47 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X24 a_2479_9004.t10 a_2479_9004.t8 a_2479_9004.t9 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X25 a_2479_9004.t18 VN.t2 a_2995_7336.t16 VSS.t43 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X26 VSS.t29 a_2080_2896.t13 a_4920_2896.t18 VSS.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X27 VOUT.t14 a_2479_7336.t23 VDD.t69 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X28 VSS.t122 VSS.t121 VSS.t122 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X29 VDD.t51 VDD.t49 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X30 a_2995_7336.t13 VP.t1 a_2479_7336.t3 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X31 VSS.t120 VSS.t119 VSS.t120 VSS.t60 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X32 a_3758_2896.t11 a_2080_2896.t14 VSS.t42 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X33 a_4920_2896.t17 a_2080_2896.t15 VSS.t35 VSS.t34 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X34 a_2479_7336.t2 VP.t2 a_2995_7336.t12 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X35 a_3758_2896.t10 a_2080_2896.t16 VSS.t32 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X36 VOUT.t16 a_2479_7336.t24 VDD.t68 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X37 VSS.t138 a_2080_2896.t17 a_3758_2896.t9 VSS.t53 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X38 a_4920_2896.t26 a_4920_2896.t25 a_4920_2896.t26 VSS.t57 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X39 a_4920_2896.t16 a_2080_2896.t18 VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X40 a_3758_2896.t8 a_2080_2896.t19 VSS.t134 VSS.t55 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X41 a_3758_2896.t7 a_2080_2896.t20 VSS.t136 VSS.t91 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X42 a_4920_2896.t24 EN.t0 VOUT.t0 VSS.t18 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X43 a_2995_7336.t11 VP.t3 a_2479_7336.t15 VSS.t60 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X44 VDD.t8 a_2479_9004.t6 a_2479_9004.t7 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X45 VOUT.t13 VOUT.t11 VOUT.t12 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X46 a_4920_2896.t15 a_2080_2896.t21 VSS.t137 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X47 VDD.t48 VDD.t47 VDD.t48 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X48 VSS.t44 a_2080_2896.t22 a_4920_2896.t14 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X49 VDD.t46 VDD.t45 VDD.t46 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X50 VSS.t118 VSS.t117 VSS.t118 VSS.t33 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X51 VDD.t67 a_2479_7336.t25 VOUT.t27 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X52 VSS.t116 VSS.t114 VSS.t115 VSS.t77 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X53 VSS.t113 VSS.t112 VSS.t113 VSS.t60 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X54 VOUT.t10 VOUT.t8 VOUT.t9 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X55 VSS.t46 a_2080_2896.t23 a_4920_2896.t13 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X56 VOUT.t7 VOUT.t6 VOUT.t7 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X57 a_2995_7336.t15 VN.t3 a_2479_9004.t17 VSS.t60 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X58 VDD.t66 a_2479_7336.t26 VOUT.t23 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X59 VSS.t111 VSS.t109 VSS.t110 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X60 VDD.t44 VDD.t42 VDD.t43 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X61 a_2479_9004.t5 a_2479_9004.t4 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X62 C1.t1 VOUT.t1 sky130_fd_pr__cap_mim_m3_1 l=25.5 w=25.5
X63 VDD.t65 a_2479_7336.t27 VOUT.t22 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X64 VSS.t133 a_2080_2896.t24 a_3758_2896.t6 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X65 a_4920_2896.t12 a_2080_2896.t25 VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X66 VSS.t108 VSS.t107 VSS.t108 VSS.t33 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X67 VOUT.t30 a_2479_7336.t28 VDD.t64 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X68 VDD.t76 a_2479_9004.t21 a_2479_7336.t17 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X69 VDD.t41 VDD.t40 VDD.t41 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X70 VSS.t106 VSS.t105 VSS.t106 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X71 VDD.t39 VDD.t38 VDD.t39 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X72 VOUT.t29 a_2479_7336.t29 VDD.t63 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X73 VSS.t1 a_2080_2896.t26 a_3758_2896.t5 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X74 VSS.t104 VSS.t103 VSS.t104 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X75 VDD.t37 VDD.t36 VDD.t37 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X76 VSS.t102 VSS.t101 VSS.t102 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X77 VDD.t35 VDD.t33 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X78 a_3758_2896.t4 a_2080_2896.t27 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X79 VSS.t100 VSS.t99 VSS.t100 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X80 VSS.t98 VSS.t97 VSS.t98 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X81 VSS.t96 VSS.t95 VSS.t96 VSS.t88 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X82 a_2995_7336.t10 VP.t4 a_2479_7336.t16 VSS.t33 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X83 VSS.t94 VSS.t93 VSS.t94 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X84 a_4920_2896.t11 a_2080_2896.t28 VSS.t28 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X85 a_2479_7336.t6 VP.t5 a_2995_7336.t9 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X86 a_2080_2896.t2 a_2080_2896.t0 a_2080_2896.t1 VSS.t59 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X87 a_2479_7336.t1 a_2479_9004.t22 VDD.t4 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X88 VSS.t51 a_2080_2896.t29 a_4920_2896.t10 VSS.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X89 a_2995_7336.t0 VN.t4 a_2479_9004.t16 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X90 VOUT.t28 a_2479_7336.t30 VDD.t62 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X91 a_4920_2896.t9 a_2080_2896.t30 VSS.t50 VSS.t34 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X92 a_2479_9004.t15 VN.t5 a_2995_7336.t4 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X93 VDD.t56 a_2479_9004.t23 a_2479_7336.t9 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X94 VDD.t32 VDD.t30 VDD.t32 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X95 VSS.t62 a_2080_2896.t31 a_4920_2896.t8 VSS.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X96 VOUT.t17 a_2479_7336.t31 VDD.t61 VDD.t50 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X97 VSS.t63 a_2080_2896.t32 a_4920_2896.t7 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X98 a_2995_7336.t5 VN.t6 a_2479_9004.t14 VSS.t33 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X99 VDD.t29 VDD.t27 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X100 a_4920_2896.t6 a_2080_2896.t33 VSS.t54 VSS.t53 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X101 a_2479_9004.t13 VN.t7 a_2995_7336.t3 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X102 VSS.t61 a_2080_2896.t34 a_4920_2896.t5 VSS.t55 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X103 VSS.t92 VSS.t90 VSS.t92 VSS.t91 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X104 a_2995_7336.t8 VP.t6 a_2479_7336.t5 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X105 a_2479_7336.t4 VP.t7 a_2995_7336.t7 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X106 VSS.t89 VSS.t87 VSS.t89 VSS.t88 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X107 VSS.t37 a_2080_2896.t35 a_3758_2896.t3 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X108 VSS.t4 a_2080_2896.t36 a_3758_2896.t2 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X109 VSS.t86 VSS.t84 VSS.t85 VSS.t77 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X110 a_3758_2896.t1 a_2080_2896.t37 VSS.t25 VSS.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X111 VDD.t6 a_2479_9004.t2 a_2479_9004.t3 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X112 VSS.t45 a_2080_2896.t38 a_3758_2896.t0 VSS.t34 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X113 IBIAS.t1 IBIAS.t0 IBIAS.t1 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X114 VSS.t83 VSS.t82 VSS.t83 VSS.t43 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X115 VDD.t26 VDD.t25 VDD.t26 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X116 VSS.t27 a_2080_2896.t39 a_4920_2896.t4 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X117 VDD.t24 VDD.t22 VDD.t23 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X118 IBIAS.t2 EN.t1 a_2080_2896.t7 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X119 VSS.t81 VSS.t80 VSS.t81 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X120 a_2479_7336.t0 a_2479_9004.t24 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X121 a_4920_2896.t3 a_2080_2896.t40 VSS.t48 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X122 a_4920_2896.t2 a_2080_2896.t41 VSS.t40 VSS.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X123 VOUT.t31 a_2479_7336.t32 VDD.t60 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X124 a_2479_7336.t8 C1.t0 VSS.t49 sky130_fd_pr__res_xhigh_po_1p41 l=14
X125 VDD.t21 VDD.t19 VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X126 VDD.t18 VDD.t16 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X127 a_3758_2896.t14 a_3758_2896.t13 a_3758_2896.t14 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X128 VOUT.t19 a_2479_7336.t33 VDD.t59 VDD.t7 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X129 VOUT.t5 VOUT.t4 VOUT.t5 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X130 a_4920_2896.t1 a_2080_2896.t42 VSS.t135 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X131 a_3758_2896.t12 EN.t2 a_2995_7336.t1 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X132 VSS.t41 a_2080_2896.t43 a_4920_2896.t0 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X133 VOUT.t3 VOUT.t2 VOUT.t3 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X134 VOUT.t20 a_2479_7336.t34 VDD.t58 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X135 VSS.t79 VSS.t76 VSS.t78 VSS.t77 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X136 a_2995_7336.t19 a_2995_7336.t17 a_2995_7336.t18 VSS.t52 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X137 VDD.t15 VDD.t13 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X138 VSS.t75 VSS.t74 VSS.t75 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X139 VDD.t12 VDD.t9 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X140 a_2080_2896.t4 a_2080_2896.t3 VSS.t31 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X141 VSS.t73 VSS.t71 VSS.t72 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X142 VSS.t70 VSS.t69 VSS.t70 VSS.t43 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X143 VDD.t57 a_2479_7336.t35 VOUT.t21 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X144 VSS.t68 VSS.t67 VSS.t68 VSS.t30 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X145 a_2479_9004.t1 a_2479_9004.t0 VDD.t75 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X146 VSS.t66 VSS.t65 VSS.t66 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
R0 VSS.n2312 VSS.n144 2542.66
R1 VSS.n2145 VSS.n2134 1321.06
R2 VSS.n2147 VSS.n2132 1321.06
R3 VSS.n2314 VSS.n140 1321.06
R4 VSS.n2307 VSS.n2306 1321.06
R5 VSS.n1540 VSS.n636 1268.91
R6 VSS.n2622 VSS.n37 1268.91
R7 VSS.n1496 VSS.n1495 1268.91
R8 VSS.n2594 VSS.n41 1268.91
R9 VSS.n1627 VSS.n572 1268.91
R10 VSS.n1595 VSS.n604 1268.91
R11 VSS.n987 VSS.n570 1268.91
R12 VSS.n1552 VSS.n1551 1268.91
R13 VSS.n1343 VSS.n1279 1268.91
R14 VSS.n1643 VSS.n509 1268.91
R15 VSS.n1302 VSS.n1276 1268.91
R16 VSS.n1645 VSS.n506 1268.91
R17 VSS.n1829 VSS.n375 1182
R18 VSS.n2003 VSS.n342 1182
R19 VSS.n1832 VSS.n377 1182
R20 VSS.n1921 VSS.n340 1182
R21 VSS.n1093 VSS.n1091 1182
R22 VSS.n2396 VSS.n116 1182
R23 VSS.n2548 VSS.n2545 1182
R24 VSS.n1347 VSS.n719 1182
R25 VSS.n2406 VSS.n101 996.588
R26 VSS.n2312 VSS.n142 614.067
R27 VSS.n2454 VSS.n89 602.588
R28 VSS.n2502 VSS.n77 602.588
R29 VSS.n197 VSS.n196 585
R30 VSS.n199 VSS.n197 585
R31 VSS.n2224 VSS.n2223 585
R32 VSS.n2225 VSS.n2224 585
R33 VSS.n2222 VSS.n204 585
R34 VSS.n204 VSS.n203 585
R35 VSS.n2221 VSS.n2220 585
R36 VSS.n2220 VSS.n2219 585
R37 VSS.n206 VSS.n205 585
R38 VSS.n207 VSS.n206 585
R39 VSS.n2212 VSS.n2211 585
R40 VSS.n2213 VSS.n2212 585
R41 VSS.n2210 VSS.n212 585
R42 VSS.n212 VSS.n211 585
R43 VSS.n2209 VSS.n2208 585
R44 VSS.n2208 VSS.n2207 585
R45 VSS.n214 VSS.n213 585
R46 VSS.n215 VSS.n214 585
R47 VSS.n2200 VSS.n2199 585
R48 VSS.n2201 VSS.n2200 585
R49 VSS.n2198 VSS.n220 585
R50 VSS.n220 VSS.n219 585
R51 VSS.n2197 VSS.n2196 585
R52 VSS.n2196 VSS.n2195 585
R53 VSS.n222 VSS.n221 585
R54 VSS.n223 VSS.n222 585
R55 VSS.n2188 VSS.n2187 585
R56 VSS.n2189 VSS.n2188 585
R57 VSS.n2186 VSS.n228 585
R58 VSS.n228 VSS.n227 585
R59 VSS.n2185 VSS.n2184 585
R60 VSS.n2184 VSS.n2183 585
R61 VSS.n230 VSS.n229 585
R62 VSS.n231 VSS.n230 585
R63 VSS.n2176 VSS.n2175 585
R64 VSS.n2177 VSS.n2176 585
R65 VSS.n2174 VSS.n236 585
R66 VSS.n236 VSS.n235 585
R67 VSS.n2173 VSS.n2172 585
R68 VSS.n2172 VSS.n2171 585
R69 VSS.n238 VSS.n237 585
R70 VSS.n2164 VSS.n238 585
R71 VSS.n2163 VSS.n2162 585
R72 VSS.n2165 VSS.n2163 585
R73 VSS.n2161 VSS.n2122 585
R74 VSS.n2122 VSS.n2121 585
R75 VSS.n2160 VSS.n2159 585
R76 VSS.n2159 VSS.n2158 585
R77 VSS.n2124 VSS.n2123 585
R78 VSS.n2125 VSS.n2124 585
R79 VSS.n2151 VSS.n2150 585
R80 VSS.n2152 VSS.n2151 585
R81 VSS.n2149 VSS.n2130 585
R82 VSS.n2130 VSS.n2129 585
R83 VSS.n2148 VSS.n2147 585
R84 VSS.n2147 VSS.n2146 585
R85 VSS.n2132 VSS.n2131 585
R86 VSS.n2138 VSS.n2136 585
R87 VSS.n2139 VSS.n2135 585
R88 VSS.n2142 VSS.n2141 585
R89 VSS.n2143 VSS.n2134 585
R90 VSS.n2134 VSS.n2133 585
R91 VSS.n2145 VSS.n2144 585
R92 VSS.n2146 VSS.n2145 585
R93 VSS.n2128 VSS.n2127 585
R94 VSS.n2129 VSS.n2128 585
R95 VSS.n2154 VSS.n2153 585
R96 VSS.n2153 VSS.n2152 585
R97 VSS.n2155 VSS.n2126 585
R98 VSS.n2126 VSS.n2125 585
R99 VSS.n2157 VSS.n2156 585
R100 VSS.n2158 VSS.n2157 585
R101 VSS.n2120 VSS.n2119 585
R102 VSS.n2121 VSS.n2120 585
R103 VSS.n2167 VSS.n2166 585
R104 VSS.n2166 VSS.n2165 585
R105 VSS.n2168 VSS.n2118 585
R106 VSS.n2164 VSS.n2118 585
R107 VSS.n2170 VSS.n2169 585
R108 VSS.n2171 VSS.n2170 585
R109 VSS.n234 VSS.n233 585
R110 VSS.n235 VSS.n234 585
R111 VSS.n2179 VSS.n2178 585
R112 VSS.n2178 VSS.n2177 585
R113 VSS.n2180 VSS.n232 585
R114 VSS.n232 VSS.n231 585
R115 VSS.n2182 VSS.n2181 585
R116 VSS.n2183 VSS.n2182 585
R117 VSS.n226 VSS.n225 585
R118 VSS.n227 VSS.n226 585
R119 VSS.n2191 VSS.n2190 585
R120 VSS.n2190 VSS.n2189 585
R121 VSS.n2192 VSS.n224 585
R122 VSS.n224 VSS.n223 585
R123 VSS.n2194 VSS.n2193 585
R124 VSS.n2195 VSS.n2194 585
R125 VSS.n218 VSS.n217 585
R126 VSS.n219 VSS.n218 585
R127 VSS.n2203 VSS.n2202 585
R128 VSS.n2202 VSS.n2201 585
R129 VSS.n2204 VSS.n216 585
R130 VSS.n216 VSS.n215 585
R131 VSS.n2206 VSS.n2205 585
R132 VSS.n2207 VSS.n2206 585
R133 VSS.n210 VSS.n209 585
R134 VSS.n211 VSS.n210 585
R135 VSS.n2215 VSS.n2214 585
R136 VSS.n2214 VSS.n2213 585
R137 VSS.n2216 VSS.n208 585
R138 VSS.n208 VSS.n207 585
R139 VSS.n2218 VSS.n2217 585
R140 VSS.n2219 VSS.n2218 585
R141 VSS.n202 VSS.n201 585
R142 VSS.n203 VSS.n202 585
R143 VSS.n2227 VSS.n2226 585
R144 VSS.n2226 VSS.n2225 585
R145 VSS.n2228 VSS.n200 585
R146 VSS.n200 VSS.n199 585
R147 VSS.n2315 VSS.n2314 585
R148 VSS.n146 VSS.n141 585
R149 VSS.n2311 VSS.n2310 585
R150 VSS.n2312 VSS.n2311 585
R151 VSS.n2309 VSS.n145 585
R152 VSS.n2308 VSS.n2307 585
R153 VSS.n2306 VSS.n147 585
R154 VSS.n2306 VSS.n142 585
R155 VSS.n2305 VSS.n149 585
R156 VSS.n2305 VSS.n2304 585
R157 VSS.n2295 VSS.n148 585
R158 VSS.n150 VSS.n148 585
R159 VSS.n2297 VSS.n2296 585
R160 VSS.n2298 VSS.n2297 585
R161 VSS.n2294 VSS.n155 585
R162 VSS.n155 VSS.n154 585
R163 VSS.n2293 VSS.n2292 585
R164 VSS.n2292 VSS.n2291 585
R165 VSS.n157 VSS.n156 585
R166 VSS.n158 VSS.n157 585
R167 VSS.n2284 VSS.n2283 585
R168 VSS.n2285 VSS.n2284 585
R169 VSS.n2282 VSS.n163 585
R170 VSS.n163 VSS.n162 585
R171 VSS.n2281 VSS.n2280 585
R172 VSS.n2280 VSS.n2279 585
R173 VSS.n165 VSS.n164 585
R174 VSS.n166 VSS.n165 585
R175 VSS.n2272 VSS.n2271 585
R176 VSS.n2273 VSS.n2272 585
R177 VSS.n2270 VSS.n171 585
R178 VSS.n171 VSS.n170 585
R179 VSS.n2269 VSS.n2268 585
R180 VSS.n2268 VSS.n2267 585
R181 VSS.n173 VSS.n172 585
R182 VSS.n174 VSS.n173 585
R183 VSS.n2260 VSS.n2259 585
R184 VSS.n2261 VSS.n2260 585
R185 VSS.n2258 VSS.n179 585
R186 VSS.n179 VSS.n178 585
R187 VSS.n2257 VSS.n2256 585
R188 VSS.n2256 VSS.n2255 585
R189 VSS.n181 VSS.n180 585
R190 VSS.n182 VSS.n181 585
R191 VSS.n2248 VSS.n2247 585
R192 VSS.n2249 VSS.n2248 585
R193 VSS.n2246 VSS.n187 585
R194 VSS.n187 VSS.n186 585
R195 VSS.n2245 VSS.n2244 585
R196 VSS.n2244 VSS.n2243 585
R197 VSS.n189 VSS.n188 585
R198 VSS.n190 VSS.n189 585
R199 VSS.n2236 VSS.n2235 585
R200 VSS.n2237 VSS.n2236 585
R201 VSS.n2234 VSS.n195 585
R202 VSS.n195 VSS.n194 585
R203 VSS.n2233 VSS.n2232 585
R204 VSS.n2232 VSS.n2231 585
R205 VSS.n2230 VSS.n2229 585
R206 VSS.n2231 VSS.n2230 585
R207 VSS.n193 VSS.n192 585
R208 VSS.n194 VSS.n193 585
R209 VSS.n2239 VSS.n2238 585
R210 VSS.n2238 VSS.n2237 585
R211 VSS.n2240 VSS.n191 585
R212 VSS.n191 VSS.n190 585
R213 VSS.n2242 VSS.n2241 585
R214 VSS.n2243 VSS.n2242 585
R215 VSS.n185 VSS.n184 585
R216 VSS.n186 VSS.n185 585
R217 VSS.n2251 VSS.n2250 585
R218 VSS.n2250 VSS.n2249 585
R219 VSS.n2252 VSS.n183 585
R220 VSS.n183 VSS.n182 585
R221 VSS.n2254 VSS.n2253 585
R222 VSS.n2255 VSS.n2254 585
R223 VSS.n177 VSS.n176 585
R224 VSS.n178 VSS.n177 585
R225 VSS.n2263 VSS.n2262 585
R226 VSS.n2262 VSS.n2261 585
R227 VSS.n2264 VSS.n175 585
R228 VSS.n175 VSS.n174 585
R229 VSS.n2266 VSS.n2265 585
R230 VSS.n2267 VSS.n2266 585
R231 VSS.n169 VSS.n168 585
R232 VSS.n170 VSS.n169 585
R233 VSS.n2275 VSS.n2274 585
R234 VSS.n2274 VSS.n2273 585
R235 VSS.n2276 VSS.n167 585
R236 VSS.n167 VSS.n166 585
R237 VSS.n2278 VSS.n2277 585
R238 VSS.n2279 VSS.n2278 585
R239 VSS.n161 VSS.n160 585
R240 VSS.n162 VSS.n161 585
R241 VSS.n2287 VSS.n2286 585
R242 VSS.n2286 VSS.n2285 585
R243 VSS.n2288 VSS.n159 585
R244 VSS.n159 VSS.n158 585
R245 VSS.n2290 VSS.n2289 585
R246 VSS.n2291 VSS.n2290 585
R247 VSS.n153 VSS.n152 585
R248 VSS.n154 VSS.n153 585
R249 VSS.n2300 VSS.n2299 585
R250 VSS.n2299 VSS.n2298 585
R251 VSS.n2301 VSS.n151 585
R252 VSS.n151 VSS.n150 585
R253 VSS.n2303 VSS.n2302 585
R254 VSS.n2304 VSS.n2303 585
R255 VSS.n140 VSS.n138 585
R256 VSS.n142 VSS.n140 585
R257 VSS.n1641 VSS.n509 585
R258 VSS.n1640 VSS.n1639 585
R259 VSS.n512 VSS.n511 585
R260 VSS.n1637 VSS.n512 585
R261 VSS.n525 VSS.n524 585
R262 VSS.n527 VSS.n526 585
R263 VSS.n529 VSS.n528 585
R264 VSS.n531 VSS.n530 585
R265 VSS.n533 VSS.n532 585
R266 VSS.n535 VSS.n534 585
R267 VSS.n537 VSS.n536 585
R268 VSS.n539 VSS.n538 585
R269 VSS.n541 VSS.n540 585
R270 VSS.n543 VSS.n542 585
R271 VSS.n545 VSS.n544 585
R272 VSS.n547 VSS.n546 585
R273 VSS.n549 VSS.n548 585
R274 VSS.n551 VSS.n550 585
R275 VSS.n553 VSS.n552 585
R276 VSS.n555 VSS.n554 585
R277 VSS.n557 VSS.n556 585
R278 VSS.n558 VSS.n523 585
R279 VSS.n561 VSS.n560 585
R280 VSS.n559 VSS.n506 585
R281 VSS.n1646 VSS.n1645 585
R282 VSS.n1645 VSS.n1644 585
R283 VSS.n505 VSS.n504 585
R284 VSS.n1378 VSS.n505 585
R285 VSS.n1375 VSS.n1374 585
R286 VSS.n1376 VSS.n1375 585
R287 VSS.n1372 VSS.n709 585
R288 VSS.n1412 VSS.n709 585
R289 VSS.n902 VSS.n710 585
R290 VSS.n903 VSS.n902 585
R291 VSS.n1368 VSS.n701 585
R292 VSS.n1418 VSS.n701 585
R293 VSS.n1367 VSS.n1366 585
R294 VSS.n1366 VSS.n1365 585
R295 VSS.n712 VSS.n711 585
R296 VSS.n1363 VSS.n712 585
R297 VSS.n1296 VSS.n1295 585
R298 VSS.n1295 VSS.n718 585
R299 VSS.n1297 VSS.n717 585
R300 VSS.n1357 VSS.n717 585
R301 VSS.n1299 VSS.n1298 585
R302 VSS.n1298 VSS.n1278 585
R303 VSS.n1300 VSS.n1276 585
R304 VSS.n1344 VSS.n1276 585
R305 VSS.n1303 VSS.n1302 585
R306 VSS.n1304 VSS.n1294 585
R307 VSS.n1306 VSS.n1305 585
R308 VSS.n1308 VSS.n1292 585
R309 VSS.n1310 VSS.n1309 585
R310 VSS.n1311 VSS.n1291 585
R311 VSS.n1313 VSS.n1312 585
R312 VSS.n1315 VSS.n1289 585
R313 VSS.n1317 VSS.n1316 585
R314 VSS.n1318 VSS.n1288 585
R315 VSS.n1320 VSS.n1319 585
R316 VSS.n1322 VSS.n1286 585
R317 VSS.n1324 VSS.n1323 585
R318 VSS.n1325 VSS.n1285 585
R319 VSS.n1327 VSS.n1326 585
R320 VSS.n1329 VSS.n1283 585
R321 VSS.n1331 VSS.n1330 585
R322 VSS.n1332 VSS.n1282 585
R323 VSS.n1334 VSS.n1333 585
R324 VSS.n1336 VSS.n1281 585
R325 VSS.n1337 VSS.n1280 585
R326 VSS.n1340 VSS.n1339 585
R327 VSS.n1341 VSS.n1279 585
R328 VSS.n1279 VSS.n723 585
R329 VSS.n1343 VSS.n1342 585
R330 VSS.n1344 VSS.n1343 585
R331 VSS.n716 VSS.n715 585
R332 VSS.n1278 VSS.n716 585
R333 VSS.n1359 VSS.n1358 585
R334 VSS.n1358 VSS.n1357 585
R335 VSS.n1360 VSS.n714 585
R336 VSS.n718 VSS.n714 585
R337 VSS.n1362 VSS.n1361 585
R338 VSS.n1363 VSS.n1362 585
R339 VSS.n705 VSS.n703 585
R340 VSS.n1365 VSS.n703 585
R341 VSS.n1417 VSS.n1416 585
R342 VSS.n1418 VSS.n1417 585
R343 VSS.n1415 VSS.n704 585
R344 VSS.n903 VSS.n704 585
R345 VSS.n1414 VSS.n1413 585
R346 VSS.n1413 VSS.n1412 585
R347 VSS.n707 VSS.n706 585
R348 VSS.n1376 VSS.n707 585
R349 VSS.n510 VSS.n508 585
R350 VSS.n1378 VSS.n508 585
R351 VSS.n1643 VSS.n1642 585
R352 VSS.n1644 VSS.n1643 585
R353 VSS.n1596 VSS.n1595 585
R354 VSS.n607 VSS.n606 585
R355 VSS.n1592 VSS.n1591 585
R356 VSS.n1593 VSS.n1592 585
R357 VSS.n1590 VSS.n619 585
R358 VSS.n1589 VSS.n1588 585
R359 VSS.n1587 VSS.n1586 585
R360 VSS.n1585 VSS.n1584 585
R361 VSS.n1583 VSS.n1582 585
R362 VSS.n1581 VSS.n1580 585
R363 VSS.n1579 VSS.n1578 585
R364 VSS.n1577 VSS.n1576 585
R365 VSS.n1575 VSS.n1574 585
R366 VSS.n1573 VSS.n1572 585
R367 VSS.n1571 VSS.n1570 585
R368 VSS.n1569 VSS.n1568 585
R369 VSS.n1567 VSS.n1566 585
R370 VSS.n1565 VSS.n1564 585
R371 VSS.n1563 VSS.n1562 585
R372 VSS.n1561 VSS.n1560 585
R373 VSS.n1559 VSS.n1558 585
R374 VSS.n1557 VSS.n1556 585
R375 VSS.n1555 VSS.n1554 585
R376 VSS.n1553 VSS.n1552 585
R377 VSS.n1551 VSS.n620 585
R378 VSS.n1551 VSS.n1550 585
R379 VSS.n999 VSS.n601 585
R380 VSS.n1600 VSS.n601 585
R381 VSS.n1050 VSS.n1000 585
R382 VSS.n1050 VSS.n1049 585
R383 VSS.n1052 VSS.n1051 585
R384 VSS.n1051 VSS.n595 585
R385 VSS.n997 VSS.n594 585
R386 VSS.n1608 VSS.n594 585
R387 VSS.n995 VSS.n994 585
R388 VSS.n994 VSS.n993 585
R389 VSS.n1057 VSS.n587 585
R390 VSS.n1614 VSS.n587 585
R391 VSS.n1060 VSS.n1059 585
R392 VSS.n1060 VSS.n586 585
R393 VSS.n1062 VSS.n1061 585
R394 VSS.n1061 VSS.n578 585
R395 VSS.n990 VSS.n577 585
R396 VSS.n1622 VSS.n577 585
R397 VSS.n1067 VSS.n1066 585
R398 VSS.n1068 VSS.n1067 585
R399 VSS.n989 VSS.n570 585
R400 VSS.n1628 VSS.n570 585
R401 VSS.n988 VSS.n987 585
R402 VSS.n985 VSS.n934 585
R403 VSS.n984 VSS.n983 585
R404 VSS.n982 VSS.n981 585
R405 VSS.n980 VSS.n936 585
R406 VSS.n978 VSS.n977 585
R407 VSS.n976 VSS.n937 585
R408 VSS.n975 VSS.n974 585
R409 VSS.n972 VSS.n938 585
R410 VSS.n970 VSS.n969 585
R411 VSS.n968 VSS.n939 585
R412 VSS.n967 VSS.n966 585
R413 VSS.n964 VSS.n940 585
R414 VSS.n962 VSS.n961 585
R415 VSS.n960 VSS.n941 585
R416 VSS.n959 VSS.n958 585
R417 VSS.n956 VSS.n942 585
R418 VSS.n954 VSS.n953 585
R419 VSS.n952 VSS.n943 585
R420 VSS.n951 VSS.n950 585
R421 VSS.n948 VSS.n944 585
R422 VSS.n946 VSS.n945 585
R423 VSS.n574 VSS.n572 585
R424 VSS.n572 VSS.n569 585
R425 VSS.n1627 VSS.n1626 585
R426 VSS.n1628 VSS.n1627 585
R427 VSS.n1625 VSS.n573 585
R428 VSS.n1068 VSS.n573 585
R429 VSS.n1624 VSS.n1623 585
R430 VSS.n1623 VSS.n1622 585
R431 VSS.n576 VSS.n575 585
R432 VSS.n578 VSS.n576 585
R433 VSS.n590 VSS.n588 585
R434 VSS.n588 VSS.n586 585
R435 VSS.n1613 VSS.n1612 585
R436 VSS.n1614 VSS.n1613 585
R437 VSS.n1611 VSS.n589 585
R438 VSS.n993 VSS.n589 585
R439 VSS.n1610 VSS.n1609 585
R440 VSS.n1609 VSS.n1608 585
R441 VSS.n592 VSS.n591 585
R442 VSS.n595 VSS.n592 585
R443 VSS.n605 VSS.n603 585
R444 VSS.n1049 VSS.n603 585
R445 VSS.n1599 VSS.n1598 585
R446 VSS.n1600 VSS.n1599 585
R447 VSS.n1597 VSS.n604 585
R448 VSS.n1550 VSS.n604 585
R449 VSS.n2622 VSS.n2621 585
R450 VSS.n2620 VSS.n36 585
R451 VSS.n2619 VSS.n35 585
R452 VSS.n2624 VSS.n35 585
R453 VSS.n2618 VSS.n2617 585
R454 VSS.n2616 VSS.n2615 585
R455 VSS.n2614 VSS.n2613 585
R456 VSS.n2612 VSS.n2611 585
R457 VSS.n2610 VSS.n2609 585
R458 VSS.n2607 VSS.n2606 585
R459 VSS.n2605 VSS.n2604 585
R460 VSS.n27 VSS.n26 585
R461 VSS.n29 VSS.n28 585
R462 VSS.n19 VSS.n18 585
R463 VSS.n2627 VSS.n2626 585
R464 VSS.n2579 VSS.n20 585
R465 VSS.n2581 VSS.n2580 585
R466 VSS.n2583 VSS.n2582 585
R467 VSS.n2585 VSS.n2584 585
R468 VSS.n2587 VSS.n2586 585
R469 VSS.n2589 VSS.n2588 585
R470 VSS.n2591 VSS.n2590 585
R471 VSS.n2593 VSS.n2592 585
R472 VSS.n2595 VSS.n2594 585
R473 VSS.n2596 VSS.n41 585
R474 VSS.n41 VSS.n21 585
R475 VSS.n2598 VSS.n2597 585
R476 VSS.n2599 VSS.n2598 585
R477 VSS.n2578 VSS.n40 585
R478 VSS.n45 VSS.n40 585
R479 VSS.n2577 VSS.n2576 585
R480 VSS.n2576 VSS.n2575 585
R481 VSS.n43 VSS.n42 585
R482 VSS.n44 VSS.n43 585
R483 VSS.n2568 VSS.n2567 585
R484 VSS.n2569 VSS.n2568 585
R485 VSS.n2566 VSS.n49 585
R486 VSS.n2546 VSS.n49 585
R487 VSS.n2565 VSS.n2564 585
R488 VSS.n2564 VSS.n2563 585
R489 VSS.n51 VSS.n50 585
R490 VSS.n57 VSS.n51 585
R491 VSS.n640 VSS.n56 585
R492 VSS.n2557 VSS.n56 585
R493 VSS.n642 VSS.n641 585
R494 VSS.n644 VSS.n642 585
R495 VSS.n1495 VSS.n639 585
R496 VSS.n1495 VSS.n1494 585
R497 VSS.n1497 VSS.n1496 585
R498 VSS.n1499 VSS.n1498 585
R499 VSS.n1501 VSS.n1500 585
R500 VSS.n1503 VSS.n1502 585
R501 VSS.n1505 VSS.n1504 585
R502 VSS.n1507 VSS.n1506 585
R503 VSS.n1509 VSS.n1508 585
R504 VSS.n1511 VSS.n1510 585
R505 VSS.n1513 VSS.n1512 585
R506 VSS.n1515 VSS.n1514 585
R507 VSS.n1517 VSS.n1516 585
R508 VSS.n1519 VSS.n1518 585
R509 VSS.n1521 VSS.n1520 585
R510 VSS.n1523 VSS.n1522 585
R511 VSS.n1525 VSS.n1524 585
R512 VSS.n1527 VSS.n1526 585
R513 VSS.n1529 VSS.n1528 585
R514 VSS.n1531 VSS.n1530 585
R515 VSS.n1533 VSS.n1532 585
R516 VSS.n1535 VSS.n1534 585
R517 VSS.n1537 VSS.n1536 585
R518 VSS.n1538 VSS.n637 585
R519 VSS.n1540 VSS.n1539 585
R520 VSS.n1541 VSS.n1540 585
R521 VSS.n638 VSS.n636 585
R522 VSS.n1494 VSS.n636 585
R523 VSS.n55 VSS.n54 585
R524 VSS.n644 VSS.n55 585
R525 VSS.n2559 VSS.n2558 585
R526 VSS.n2558 VSS.n2557 585
R527 VSS.n2560 VSS.n53 585
R528 VSS.n57 VSS.n53 585
R529 VSS.n2562 VSS.n2561 585
R530 VSS.n2563 VSS.n2562 585
R531 VSS.n48 VSS.n47 585
R532 VSS.n2546 VSS.n48 585
R533 VSS.n2571 VSS.n2570 585
R534 VSS.n2570 VSS.n2569 585
R535 VSS.n2572 VSS.n46 585
R536 VSS.n46 VSS.n44 585
R537 VSS.n2574 VSS.n2573 585
R538 VSS.n2575 VSS.n2574 585
R539 VSS.n39 VSS.n38 585
R540 VSS.n45 VSS.n39 585
R541 VSS.n2601 VSS.n2600 585
R542 VSS.n2600 VSS.n2599 585
R543 VSS.n2602 VSS.n37 585
R544 VSS.n37 VSS.n21 585
R545 VSS.n2001 VSS.n342 585
R546 VSS.n2000 VSS.n1999 585
R547 VSS.n1997 VSS.n343 585
R548 VSS.n1997 VSS.n341 585
R549 VSS.n1996 VSS.n1995 585
R550 VSS.n1994 VSS.n1993 585
R551 VSS.n1992 VSS.n345 585
R552 VSS.n1990 VSS.n1989 585
R553 VSS.n1988 VSS.n346 585
R554 VSS.n1987 VSS.n1986 585
R555 VSS.n1984 VSS.n347 585
R556 VSS.n1982 VSS.n1981 585
R557 VSS.n1980 VSS.n348 585
R558 VSS.n1979 VSS.n1978 585
R559 VSS.n1976 VSS.n349 585
R560 VSS.n1974 VSS.n1973 585
R561 VSS.n351 VSS.n350 585
R562 VSS.n1969 VSS.n1968 585
R563 VSS.n1966 VSS.n1965 585
R564 VSS.n1964 VSS.n1963 585
R565 VSS.n1962 VSS.n1961 585
R566 VSS.n1952 VSS.n357 585
R567 VSS.n1953 VSS.n360 585
R568 VSS.n1956 VSS.n1955 585
R569 VSS.n1951 VSS.n1950 585
R570 VSS.n1949 VSS.n1948 585
R571 VSS.n1947 VSS.n364 585
R572 VSS.n1945 VSS.n1944 585
R573 VSS.n1943 VSS.n365 585
R574 VSS.n1942 VSS.n1941 585
R575 VSS.n1939 VSS.n366 585
R576 VSS.n1937 VSS.n1936 585
R577 VSS.n1935 VSS.n367 585
R578 VSS.n1934 VSS.n1933 585
R579 VSS.n1931 VSS.n368 585
R580 VSS.n1929 VSS.n1928 585
R581 VSS.n1927 VSS.n369 585
R582 VSS.n1926 VSS.n1925 585
R583 VSS.n1923 VSS.n370 585
R584 VSS.n1921 VSS.n1920 585
R585 VSS.n1919 VSS.n340 585
R586 VSS.n2004 VSS.n340 585
R587 VSS.n1918 VSS.n339 585
R588 VSS.n2005 VSS.n339 585
R589 VSS.n1917 VSS.n338 585
R590 VSS.n2006 VSS.n338 585
R591 VSS.n1916 VSS.n1915 585
R592 VSS.n1915 VSS.n334 585
R593 VSS.n1914 VSS.n333 585
R594 VSS.n2012 VSS.n333 585
R595 VSS.n1913 VSS.n332 585
R596 VSS.n2013 VSS.n332 585
R597 VSS.n1912 VSS.n331 585
R598 VSS.n2014 VSS.n331 585
R599 VSS.n1911 VSS.n1910 585
R600 VSS.n1910 VSS.n327 585
R601 VSS.n1909 VSS.n326 585
R602 VSS.n2020 VSS.n326 585
R603 VSS.n1908 VSS.n325 585
R604 VSS.n2021 VSS.n325 585
R605 VSS.n1907 VSS.n324 585
R606 VSS.n2022 VSS.n324 585
R607 VSS.n1906 VSS.n1905 585
R608 VSS.n1905 VSS.n320 585
R609 VSS.n1904 VSS.n319 585
R610 VSS.n2028 VSS.n319 585
R611 VSS.n1903 VSS.n318 585
R612 VSS.n2029 VSS.n318 585
R613 VSS.n1902 VSS.n317 585
R614 VSS.n2030 VSS.n317 585
R615 VSS.n1901 VSS.n1900 585
R616 VSS.n1900 VSS.n313 585
R617 VSS.n1899 VSS.n312 585
R618 VSS.n2036 VSS.n312 585
R619 VSS.n1898 VSS.n311 585
R620 VSS.n2037 VSS.n311 585
R621 VSS.n1897 VSS.n310 585
R622 VSS.n2038 VSS.n310 585
R623 VSS.n1896 VSS.n1895 585
R624 VSS.n1895 VSS.n306 585
R625 VSS.n1894 VSS.n305 585
R626 VSS.n2044 VSS.n305 585
R627 VSS.n1893 VSS.n304 585
R628 VSS.n2045 VSS.n304 585
R629 VSS.n1892 VSS.n303 585
R630 VSS.n2046 VSS.n303 585
R631 VSS.n1891 VSS.n1890 585
R632 VSS.n1890 VSS.n299 585
R633 VSS.n1889 VSS.n298 585
R634 VSS.n2052 VSS.n298 585
R635 VSS.n1888 VSS.n297 585
R636 VSS.n2053 VSS.n297 585
R637 VSS.n1887 VSS.n296 585
R638 VSS.n2054 VSS.n296 585
R639 VSS.n1886 VSS.n1885 585
R640 VSS.n1885 VSS.n292 585
R641 VSS.n1884 VSS.n291 585
R642 VSS.n2060 VSS.n291 585
R643 VSS.n1883 VSS.n290 585
R644 VSS.n2061 VSS.n290 585
R645 VSS.n1882 VSS.n289 585
R646 VSS.n2062 VSS.n289 585
R647 VSS.n1881 VSS.n1880 585
R648 VSS.n1880 VSS.n285 585
R649 VSS.n1879 VSS.n284 585
R650 VSS.n2068 VSS.n284 585
R651 VSS.n1878 VSS.n283 585
R652 VSS.n2069 VSS.n283 585
R653 VSS.n1877 VSS.n282 585
R654 VSS.n2070 VSS.n282 585
R655 VSS.n1876 VSS.n1875 585
R656 VSS.n1875 VSS.n278 585
R657 VSS.n1874 VSS.n277 585
R658 VSS.n2076 VSS.n277 585
R659 VSS.n1873 VSS.n276 585
R660 VSS.n2077 VSS.n276 585
R661 VSS.n1872 VSS.n275 585
R662 VSS.n2078 VSS.n275 585
R663 VSS.n1871 VSS.n1870 585
R664 VSS.n1870 VSS.n274 585
R665 VSS.n1869 VSS.n270 585
R666 VSS.n2084 VSS.n270 585
R667 VSS.n1868 VSS.n269 585
R668 VSS.n2085 VSS.n269 585
R669 VSS.n1867 VSS.n268 585
R670 VSS.n2086 VSS.n268 585
R671 VSS.n1866 VSS.n1865 585
R672 VSS.n1865 VSS.n267 585
R673 VSS.n1864 VSS.n263 585
R674 VSS.n2092 VSS.n263 585
R675 VSS.n1863 VSS.n262 585
R676 VSS.n2093 VSS.n262 585
R677 VSS.n1862 VSS.n261 585
R678 VSS.n2094 VSS.n261 585
R679 VSS.n1861 VSS.n1860 585
R680 VSS.n1860 VSS.n260 585
R681 VSS.n1859 VSS.n256 585
R682 VSS.n2100 VSS.n256 585
R683 VSS.n1858 VSS.n255 585
R684 VSS.n2101 VSS.n255 585
R685 VSS.n1857 VSS.n254 585
R686 VSS.n2102 VSS.n254 585
R687 VSS.n1856 VSS.n1855 585
R688 VSS.n1855 VSS.n253 585
R689 VSS.n1854 VSS.n249 585
R690 VSS.n2108 VSS.n249 585
R691 VSS.n1853 VSS.n248 585
R692 VSS.n2109 VSS.n248 585
R693 VSS.n1852 VSS.n247 585
R694 VSS.n2110 VSS.n247 585
R695 VSS.n1851 VSS.n1850 585
R696 VSS.n1850 VSS.n246 585
R697 VSS.n1849 VSS.n240 585
R698 VSS.n2116 VSS.n240 585
R699 VSS.n1848 VSS.n1847 585
R700 VSS.n1847 VSS.n239 585
R701 VSS.n1846 VSS.n371 585
R702 VSS.n1846 VSS.n1845 585
R703 VSS.n1835 VSS.n372 585
R704 VSS.n1838 VSS.n372 585
R705 VSS.n1837 VSS.n1836 585
R706 VSS.n1839 VSS.n1837 585
R707 VSS.n1834 VSS.n377 585
R708 VSS.n377 VSS.n376 585
R709 VSS.n1833 VSS.n1832 585
R710 VSS.n379 VSS.n378 585
R711 VSS.n1755 VSS.n1754 585
R712 VSS.n1757 VSS.n1756 585
R713 VSS.n1759 VSS.n1758 585
R714 VSS.n1761 VSS.n1760 585
R715 VSS.n1763 VSS.n1762 585
R716 VSS.n1765 VSS.n1764 585
R717 VSS.n1767 VSS.n1766 585
R718 VSS.n1769 VSS.n1768 585
R719 VSS.n1771 VSS.n1770 585
R720 VSS.n1773 VSS.n1772 585
R721 VSS.n1775 VSS.n1774 585
R722 VSS.n1777 VSS.n1776 585
R723 VSS.n1779 VSS.n1778 585
R724 VSS.n1781 VSS.n1780 585
R725 VSS.n1783 VSS.n1782 585
R726 VSS.n407 VSS.n406 585
R727 VSS.n405 VSS.n403 585
R728 VSS.n1789 VSS.n1788 585
R729 VSS.n1791 VSS.n1790 585
R730 VSS.n1794 VSS.n1793 585
R731 VSS.n1792 VSS.n400 585
R732 VSS.n1800 VSS.n1799 585
R733 VSS.n1802 VSS.n1801 585
R734 VSS.n1804 VSS.n1803 585
R735 VSS.n1806 VSS.n1805 585
R736 VSS.n1808 VSS.n1807 585
R737 VSS.n1810 VSS.n1809 585
R738 VSS.n1812 VSS.n1811 585
R739 VSS.n1814 VSS.n1813 585
R740 VSS.n1816 VSS.n1815 585
R741 VSS.n1818 VSS.n1817 585
R742 VSS.n1820 VSS.n1819 585
R743 VSS.n1822 VSS.n1821 585
R744 VSS.n1824 VSS.n1823 585
R745 VSS.n1826 VSS.n1825 585
R746 VSS.n1827 VSS.n398 585
R747 VSS.n1829 VSS.n1828 585
R748 VSS.n1830 VSS.n1829 585
R749 VSS.n375 VSS.n374 585
R750 VSS.n376 VSS.n375 585
R751 VSS.n1841 VSS.n1840 585
R752 VSS.n1840 VSS.n1839 585
R753 VSS.n1842 VSS.n373 585
R754 VSS.n1838 VSS.n373 585
R755 VSS.n1844 VSS.n1843 585
R756 VSS.n1845 VSS.n1844 585
R757 VSS.n243 VSS.n241 585
R758 VSS.n241 VSS.n239 585
R759 VSS.n2115 VSS.n2114 585
R760 VSS.n2116 VSS.n2115 585
R761 VSS.n2113 VSS.n242 585
R762 VSS.n246 VSS.n242 585
R763 VSS.n2112 VSS.n2111 585
R764 VSS.n2111 VSS.n2110 585
R765 VSS.n245 VSS.n244 585
R766 VSS.n2109 VSS.n245 585
R767 VSS.n2107 VSS.n2106 585
R768 VSS.n2108 VSS.n2107 585
R769 VSS.n2105 VSS.n250 585
R770 VSS.n253 VSS.n250 585
R771 VSS.n2104 VSS.n2103 585
R772 VSS.n2103 VSS.n2102 585
R773 VSS.n252 VSS.n251 585
R774 VSS.n2101 VSS.n252 585
R775 VSS.n2099 VSS.n2098 585
R776 VSS.n2100 VSS.n2099 585
R777 VSS.n2097 VSS.n257 585
R778 VSS.n260 VSS.n257 585
R779 VSS.n2096 VSS.n2095 585
R780 VSS.n2095 VSS.n2094 585
R781 VSS.n259 VSS.n258 585
R782 VSS.n2093 VSS.n259 585
R783 VSS.n2091 VSS.n2090 585
R784 VSS.n2092 VSS.n2091 585
R785 VSS.n2089 VSS.n264 585
R786 VSS.n267 VSS.n264 585
R787 VSS.n2088 VSS.n2087 585
R788 VSS.n2087 VSS.n2086 585
R789 VSS.n266 VSS.n265 585
R790 VSS.n2085 VSS.n266 585
R791 VSS.n2083 VSS.n2082 585
R792 VSS.n2084 VSS.n2083 585
R793 VSS.n2081 VSS.n271 585
R794 VSS.n274 VSS.n271 585
R795 VSS.n2080 VSS.n2079 585
R796 VSS.n2079 VSS.n2078 585
R797 VSS.n273 VSS.n272 585
R798 VSS.n2077 VSS.n273 585
R799 VSS.n2075 VSS.n2074 585
R800 VSS.n2076 VSS.n2075 585
R801 VSS.n2073 VSS.n279 585
R802 VSS.n279 VSS.n278 585
R803 VSS.n2072 VSS.n2071 585
R804 VSS.n2071 VSS.n2070 585
R805 VSS.n281 VSS.n280 585
R806 VSS.n2069 VSS.n281 585
R807 VSS.n2067 VSS.n2066 585
R808 VSS.n2068 VSS.n2067 585
R809 VSS.n2065 VSS.n286 585
R810 VSS.n286 VSS.n285 585
R811 VSS.n2064 VSS.n2063 585
R812 VSS.n2063 VSS.n2062 585
R813 VSS.n288 VSS.n287 585
R814 VSS.n2061 VSS.n288 585
R815 VSS.n2059 VSS.n2058 585
R816 VSS.n2060 VSS.n2059 585
R817 VSS.n2057 VSS.n293 585
R818 VSS.n293 VSS.n292 585
R819 VSS.n2056 VSS.n2055 585
R820 VSS.n2055 VSS.n2054 585
R821 VSS.n295 VSS.n294 585
R822 VSS.n2053 VSS.n295 585
R823 VSS.n2051 VSS.n2050 585
R824 VSS.n2052 VSS.n2051 585
R825 VSS.n2049 VSS.n300 585
R826 VSS.n300 VSS.n299 585
R827 VSS.n2048 VSS.n2047 585
R828 VSS.n2047 VSS.n2046 585
R829 VSS.n302 VSS.n301 585
R830 VSS.n2045 VSS.n302 585
R831 VSS.n2043 VSS.n2042 585
R832 VSS.n2044 VSS.n2043 585
R833 VSS.n2041 VSS.n307 585
R834 VSS.n307 VSS.n306 585
R835 VSS.n2040 VSS.n2039 585
R836 VSS.n2039 VSS.n2038 585
R837 VSS.n309 VSS.n308 585
R838 VSS.n2037 VSS.n309 585
R839 VSS.n2035 VSS.n2034 585
R840 VSS.n2036 VSS.n2035 585
R841 VSS.n2033 VSS.n314 585
R842 VSS.n314 VSS.n313 585
R843 VSS.n2032 VSS.n2031 585
R844 VSS.n2031 VSS.n2030 585
R845 VSS.n316 VSS.n315 585
R846 VSS.n2029 VSS.n316 585
R847 VSS.n2027 VSS.n2026 585
R848 VSS.n2028 VSS.n2027 585
R849 VSS.n2025 VSS.n321 585
R850 VSS.n321 VSS.n320 585
R851 VSS.n2024 VSS.n2023 585
R852 VSS.n2023 VSS.n2022 585
R853 VSS.n323 VSS.n322 585
R854 VSS.n2021 VSS.n323 585
R855 VSS.n2019 VSS.n2018 585
R856 VSS.n2020 VSS.n2019 585
R857 VSS.n2017 VSS.n328 585
R858 VSS.n328 VSS.n327 585
R859 VSS.n2016 VSS.n2015 585
R860 VSS.n2015 VSS.n2014 585
R861 VSS.n330 VSS.n329 585
R862 VSS.n2013 VSS.n330 585
R863 VSS.n2011 VSS.n2010 585
R864 VSS.n2012 VSS.n2011 585
R865 VSS.n2009 VSS.n335 585
R866 VSS.n335 VSS.n334 585
R867 VSS.n2008 VSS.n2007 585
R868 VSS.n2007 VSS.n2006 585
R869 VSS.n337 VSS.n336 585
R870 VSS.n2005 VSS.n337 585
R871 VSS.n2003 VSS.n2002 585
R872 VSS.n2004 VSS.n2003 585
R873 VSS.n1348 VSS.n1347 585
R874 VSS.n722 VSS.n721 585
R875 VSS.n1274 VSS.n1273 585
R876 VSS.n1272 VSS.n759 585
R877 VSS.n1271 VSS.n1270 585
R878 VSS.n1269 VSS.n1268 585
R879 VSS.n1267 VSS.n1266 585
R880 VSS.n1265 VSS.n1264 585
R881 VSS.n1263 VSS.n1262 585
R882 VSS.n1261 VSS.n1260 585
R883 VSS.n1259 VSS.n1258 585
R884 VSS.n1257 VSS.n1256 585
R885 VSS.n1255 VSS.n1254 585
R886 VSS.n1253 VSS.n1252 585
R887 VSS.n1251 VSS.n1250 585
R888 VSS.n1249 VSS.n1248 585
R889 VSS.n1247 VSS.n1246 585
R890 VSS.n1245 VSS.n1244 585
R891 VSS.n1243 VSS.n1242 585
R892 VSS.n1241 VSS.n1240 585
R893 VSS.n1239 VSS.n1238 585
R894 VSS.n1237 VSS.n1236 585
R895 VSS.n1235 VSS.n1234 585
R896 VSS.n1233 VSS.n1232 585
R897 VSS.n1231 VSS.n1230 585
R898 VSS.n1229 VSS.n1228 585
R899 VSS.n1227 VSS.n1226 585
R900 VSS.n1225 VSS.n1224 585
R901 VSS.n1223 VSS.n1222 585
R902 VSS.n1221 VSS.n1220 585
R903 VSS.n1219 VSS.n1218 585
R904 VSS.n1217 VSS.n1216 585
R905 VSS.n1215 VSS.n1214 585
R906 VSS.n1213 VSS.n1212 585
R907 VSS.n1211 VSS.n1210 585
R908 VSS.n1209 VSS.n1208 585
R909 VSS.n1207 VSS.n1206 585
R910 VSS.n1205 VSS.n1204 585
R911 VSS.n1203 VSS.n1202 585
R912 VSS.n1201 VSS.n1200 585
R913 VSS.n1199 VSS.n1198 585
R914 VSS.n1197 VSS.n1196 585
R915 VSS.n1195 VSS.n1194 585
R916 VSS.n1193 VSS.n1192 585
R917 VSS.n1191 VSS.n1190 585
R918 VSS.n1189 VSS.n1188 585
R919 VSS.n1187 VSS.n1186 585
R920 VSS.n1185 VSS.n1184 585
R921 VSS.n1183 VSS.n1182 585
R922 VSS.n1181 VSS.n1180 585
R923 VSS.n1179 VSS.n1178 585
R924 VSS.n1177 VSS.n1176 585
R925 VSS.n1175 VSS.n1174 585
R926 VSS.n1173 VSS.n1172 585
R927 VSS.n1171 VSS.n1170 585
R928 VSS.n1169 VSS.n1168 585
R929 VSS.n1167 VSS.n1166 585
R930 VSS.n1165 VSS.n1164 585
R931 VSS.n1163 VSS.n1162 585
R932 VSS.n1161 VSS.n1160 585
R933 VSS.n1159 VSS.n1158 585
R934 VSS.n1157 VSS.n1156 585
R935 VSS.n1155 VSS.n1154 585
R936 VSS.n1153 VSS.n1152 585
R937 VSS.n1151 VSS.n1150 585
R938 VSS.n1149 VSS.n1148 585
R939 VSS.n1147 VSS.n1146 585
R940 VSS.n1145 VSS.n1144 585
R941 VSS.n1143 VSS.n1142 585
R942 VSS.n1141 VSS.n1140 585
R943 VSS.n1139 VSS.n1138 585
R944 VSS.n1137 VSS.n1136 585
R945 VSS.n1135 VSS.n1134 585
R946 VSS.n1133 VSS.n1132 585
R947 VSS.n1131 VSS.n760 585
R948 VSS.n1129 VSS.n1128 585
R949 VSS.n1127 VSS.n761 585
R950 VSS.n1126 VSS.n1125 585
R951 VSS.n1123 VSS.n762 585
R952 VSS.n1121 VSS.n1120 585
R953 VSS.n1119 VSS.n763 585
R954 VSS.n1118 VSS.n1117 585
R955 VSS.n1115 VSS.n764 585
R956 VSS.n1113 VSS.n1112 585
R957 VSS.n1111 VSS.n765 585
R958 VSS.n1110 VSS.n1109 585
R959 VSS.n1107 VSS.n766 585
R960 VSS.n1105 VSS.n1104 585
R961 VSS.n1103 VSS.n767 585
R962 VSS.n1102 VSS.n1101 585
R963 VSS.n1099 VSS.n768 585
R964 VSS.n1097 VSS.n1096 585
R965 VSS.n1095 VSS.n769 585
R966 VSS.n1094 VSS.n1093 585
R967 VSS.n1091 VSS.n770 585
R968 VSS.n1091 VSS.n1090 585
R969 VSS.n777 VSS.n771 585
R970 VSS.n1089 VSS.n771 585
R971 VSS.n1087 VSS.n1086 585
R972 VSS.n1088 VSS.n1087 585
R973 VSS.n1085 VSS.n773 585
R974 VSS.n773 VSS.n772 585
R975 VSS.n900 VSS.n775 585
R976 VSS.n901 VSS.n900 585
R977 VSS.n906 VSS.n905 585
R978 VSS.n905 VSS.n904 585
R979 VSS.n898 VSS.n897 585
R980 VSS.n897 VSS.n896 585
R981 VSS.n911 VSS.n910 585
R982 VSS.n912 VSS.n911 585
R983 VSS.n899 VSS.n895 585
R984 VSS.n913 VSS.n895 585
R985 VSS.n915 VSS.n894 585
R986 VSS.n915 VSS.n914 585
R987 VSS.n918 VSS.n917 585
R988 VSS.n917 VSS.n916 585
R989 VSS.n919 VSS.n893 585
R990 VSS.n893 VSS.n892 585
R991 VSS.n921 VSS.n920 585
R992 VSS.n922 VSS.n921 585
R993 VSS.n891 VSS.n890 585
R994 VSS.n923 VSS.n891 585
R995 VSS.n926 VSS.n925 585
R996 VSS.n925 VSS.n924 585
R997 VSS.n927 VSS.n888 585
R998 VSS.n888 VSS.n887 585
R999 VSS.n932 VSS.n931 585
R1000 VSS.n933 VSS.n932 585
R1001 VSS.n929 VSS.n889 585
R1002 VSS.n889 VSS.n886 585
R1003 VSS.n884 VSS.n882 585
R1004 VSS.n1071 VSS.n884 585
R1005 VSS.n1075 VSS.n1074 585
R1006 VSS.n1074 VSS.n1073 585
R1007 VSS.n885 VSS.n883 585
R1008 VSS.n1072 VSS.n885 585
R1009 VSS.n1017 VSS.n1016 585
R1010 VSS.n1020 VSS.n1017 585
R1011 VSS.n1024 VSS.n1023 585
R1012 VSS.n1023 VSS.n1022 585
R1013 VSS.n1019 VSS.n1018 585
R1014 VSS.n1021 VSS.n1019 585
R1015 VSS.n1006 VSS.n1004 585
R1016 VSS.n1004 VSS.n1002 585
R1017 VSS.n1047 VSS.n1046 585
R1018 VSS.n1048 VSS.n1047 585
R1019 VSS.n1045 VSS.n1005 585
R1020 VSS.n1005 VSS.n1003 585
R1021 VSS.n1044 VSS.n1043 585
R1022 VSS.n1043 VSS.n1042 585
R1023 VSS.n1040 VSS.n1007 585
R1024 VSS.n1041 VSS.n1040 585
R1025 VSS.n1039 VSS.n1009 585
R1026 VSS.n1039 VSS.n1038 585
R1027 VSS.n1012 VSS.n1008 585
R1028 VSS.n1037 VSS.n1008 585
R1029 VSS.n1035 VSS.n1034 585
R1030 VSS.n1036 VSS.n1035 585
R1031 VSS.n1033 VSS.n1011 585
R1032 VSS.n1011 VSS.n1010 585
R1033 VSS.n125 VSS.n124 585
R1034 VSS.n124 VSS.n123 585
R1035 VSS.n2352 VSS.n2351 585
R1036 VSS.n2353 VSS.n2352 585
R1037 VSS.n120 VSS.n119 585
R1038 VSS.n2354 VSS.n120 585
R1039 VSS.n2357 VSS.n2356 585
R1040 VSS.n2356 VSS.n2355 585
R1041 VSS.n122 VSS.n117 585
R1042 VSS.n122 VSS.n121 585
R1043 VSS.n2361 VSS.n116 585
R1044 VSS.n116 VSS.n105 585
R1045 VSS.n2396 VSS.n2395 585
R1046 VSS.n2394 VSS.n115 585
R1047 VSS.n2393 VSS.n114 585
R1048 VSS.n2398 VSS.n114 585
R1049 VSS.n2392 VSS.n2391 585
R1050 VSS.n2390 VSS.n2389 585
R1051 VSS.n2388 VSS.n2387 585
R1052 VSS.n2386 VSS.n2385 585
R1053 VSS.n2384 VSS.n2383 585
R1054 VSS.n2382 VSS.n2381 585
R1055 VSS.n2380 VSS.n2379 585
R1056 VSS.n2378 VSS.n2377 585
R1057 VSS.n2376 VSS.n2375 585
R1058 VSS.n2374 VSS.n2373 585
R1059 VSS.n2372 VSS.n2371 585
R1060 VSS.n2370 VSS.n2369 585
R1061 VSS.n2368 VSS.n2367 585
R1062 VSS.n2366 VSS.n2365 585
R1063 VSS.n2364 VSS.n2363 585
R1064 VSS.n2362 VSS.n103 585
R1065 VSS.n2399 VSS.n104 585
R1066 VSS.n2399 VSS.n2398 585
R1067 VSS.n2400 VSS.n102 585
R1068 VSS.n2403 VSS.n2402 585
R1069 VSS.n2404 VSS.n101 585
R1070 VSS.n101 VSS.n44 585
R1071 VSS.n2406 VSS.n2405 585
R1072 VSS.n2408 VSS.n100 585
R1073 VSS.n2411 VSS.n2410 585
R1074 VSS.n2412 VSS.n99 585
R1075 VSS.n2414 VSS.n2413 585
R1076 VSS.n2416 VSS.n98 585
R1077 VSS.n2419 VSS.n2418 585
R1078 VSS.n2420 VSS.n97 585
R1079 VSS.n2422 VSS.n2421 585
R1080 VSS.n2424 VSS.n96 585
R1081 VSS.n2427 VSS.n2426 585
R1082 VSS.n2428 VSS.n95 585
R1083 VSS.n2430 VSS.n2429 585
R1084 VSS.n2432 VSS.n94 585
R1085 VSS.n2435 VSS.n2434 585
R1086 VSS.n2436 VSS.n93 585
R1087 VSS.n2438 VSS.n2437 585
R1088 VSS.n2440 VSS.n92 585
R1089 VSS.n2443 VSS.n2442 585
R1090 VSS.n2444 VSS.n91 585
R1091 VSS.n2446 VSS.n2445 585
R1092 VSS.n2448 VSS.n90 585
R1093 VSS.n2451 VSS.n2450 585
R1094 VSS.n2452 VSS.n89 585
R1095 VSS.n2454 VSS.n2453 585
R1096 VSS.n2456 VSS.n88 585
R1097 VSS.n2459 VSS.n2458 585
R1098 VSS.n2460 VSS.n87 585
R1099 VSS.n2462 VSS.n2461 585
R1100 VSS.n2464 VSS.n86 585
R1101 VSS.n2467 VSS.n2466 585
R1102 VSS.n2468 VSS.n85 585
R1103 VSS.n2470 VSS.n2469 585
R1104 VSS.n2472 VSS.n84 585
R1105 VSS.n2475 VSS.n2474 585
R1106 VSS.n2476 VSS.n83 585
R1107 VSS.n2478 VSS.n2477 585
R1108 VSS.n2480 VSS.n82 585
R1109 VSS.n2483 VSS.n2482 585
R1110 VSS.n2484 VSS.n81 585
R1111 VSS.n2486 VSS.n2485 585
R1112 VSS.n2488 VSS.n80 585
R1113 VSS.n2491 VSS.n2490 585
R1114 VSS.n2492 VSS.n79 585
R1115 VSS.n2494 VSS.n2493 585
R1116 VSS.n2496 VSS.n78 585
R1117 VSS.n2499 VSS.n2498 585
R1118 VSS.n2500 VSS.n77 585
R1119 VSS.n2502 VSS.n2501 585
R1120 VSS.n2504 VSS.n76 585
R1121 VSS.n2507 VSS.n2506 585
R1122 VSS.n2508 VSS.n75 585
R1123 VSS.n2510 VSS.n2509 585
R1124 VSS.n2512 VSS.n74 585
R1125 VSS.n2515 VSS.n2514 585
R1126 VSS.n2516 VSS.n73 585
R1127 VSS.n2518 VSS.n2517 585
R1128 VSS.n2520 VSS.n72 585
R1129 VSS.n2523 VSS.n2522 585
R1130 VSS.n2524 VSS.n71 585
R1131 VSS.n2526 VSS.n2525 585
R1132 VSS.n2528 VSS.n70 585
R1133 VSS.n2531 VSS.n2530 585
R1134 VSS.n2532 VSS.n69 585
R1135 VSS.n2534 VSS.n2533 585
R1136 VSS.n2536 VSS.n68 585
R1137 VSS.n2539 VSS.n2538 585
R1138 VSS.n2540 VSS.n67 585
R1139 VSS.n2542 VSS.n2541 585
R1140 VSS.n2544 VSS.n66 585
R1141 VSS.n2545 VSS.n64 585
R1142 VSS.n2545 VSS.n44 585
R1143 VSS.n2549 VSS.n2548 585
R1144 VSS.n2548 VSS.n2547 585
R1145 VSS.n65 VSS.n62 585
R1146 VSS.n65 VSS.n52 585
R1147 VSS.n2553 VSS.n60 585
R1148 VSS.n60 VSS.n59 585
R1149 VSS.n2555 VSS.n2554 585
R1150 VSS.n2556 VSS.n2555 585
R1151 VSS.n1490 VSS.n58 585
R1152 VSS.n643 VSS.n58 585
R1153 VSS.n1492 VSS.n1491 585
R1154 VSS.n1493 VSS.n1492 585
R1155 VSS.n647 VSS.n646 585
R1156 VSS.n646 VSS.n645 585
R1157 VSS.n649 VSS.n648 585
R1158 VSS.n648 VSS.n624 585
R1159 VSS.n623 VSS.n622 585
R1160 VSS.n1542 VSS.n623 585
R1161 VSS.n1545 VSS.n1544 585
R1162 VSS.n1544 VSS.n1543 585
R1163 VSS.n1546 VSS.n621 585
R1164 VSS.n621 VSS.n608 585
R1165 VSS.n1548 VSS.n1547 585
R1166 VSS.n1549 VSS.n1548 585
R1167 VSS.n600 VSS.n599 585
R1168 VSS.n602 VSS.n600 585
R1169 VSS.n1603 VSS.n1602 585
R1170 VSS.n1602 VSS.n1601 585
R1171 VSS.n1604 VSS.n597 585
R1172 VSS.n1001 VSS.n597 585
R1173 VSS.n1606 VSS.n1605 585
R1174 VSS.n1607 VSS.n1606 585
R1175 VSS.n1389 VSS.n596 585
R1176 VSS.n596 VSS.n593 585
R1177 VSS.n584 VSS.n583 585
R1178 VSS.n992 VSS.n584 585
R1179 VSS.n1617 VSS.n1616 585
R1180 VSS.n1616 VSS.n1615 585
R1181 VSS.n1618 VSS.n580 585
R1182 VSS.n585 VSS.n580 585
R1183 VSS.n1620 VSS.n1619 585
R1184 VSS.n1621 VSS.n1620 585
R1185 VSS.n581 VSS.n579 585
R1186 VSS.n1070 VSS.n579 585
R1187 VSS.n1398 VSS.n1397 585
R1188 VSS.n1397 VSS.n571 585
R1189 VSS.n568 VSS.n567 585
R1190 VSS.n1629 VSS.n568 585
R1191 VSS.n1632 VSS.n1631 585
R1192 VSS.n1631 VSS.n1630 585
R1193 VSS.n1633 VSS.n565 585
R1194 VSS.n565 VSS.n563 585
R1195 VSS.n1635 VSS.n1634 585
R1196 VSS.n1636 VSS.n1635 585
R1197 VSS.n566 VSS.n564 585
R1198 VSS.n564 VSS.n513 585
R1199 VSS.n1384 VSS.n1382 585
R1200 VSS.n1384 VSS.n1383 585
R1201 VSS.n1386 VSS.n1385 585
R1202 VSS.n1385 VSS.n507 585
R1203 VSS.n1387 VSS.n1380 585
R1204 VSS.n1380 VSS.n1379 585
R1205 VSS.n1410 VSS.n1409 585
R1206 VSS.n1411 VSS.n1410 585
R1207 VSS.n1381 VSS.n1377 585
R1208 VSS.n1377 VSS.n708 585
R1209 VSS.n700 VSS.n698 585
R1210 VSS.n702 VSS.n700 585
R1211 VSS.n1421 VSS.n1420 585
R1212 VSS.n1420 VSS.n1419 585
R1213 VSS.n699 VSS.n697 585
R1214 VSS.n1364 VSS.n699 585
R1215 VSS.n1351 VSS.n720 585
R1216 VSS.n720 VSS.n713 585
R1217 VSS.n1355 VSS.n1354 585
R1218 VSS.n1356 VSS.n1355 585
R1219 VSS.n1349 VSS.n719 585
R1220 VSS.n1277 VSS.n719 585
R1221 VSS.n1840 VSS.n375 394
R1222 VSS.n1840 VSS.n373 394
R1223 VSS.n1844 VSS.n373 394
R1224 VSS.n1844 VSS.n241 394
R1225 VSS.n2115 VSS.n241 394
R1226 VSS.n2115 VSS.n242 394
R1227 VSS.n2111 VSS.n242 394
R1228 VSS.n2111 VSS.n245 394
R1229 VSS.n2107 VSS.n245 394
R1230 VSS.n2107 VSS.n250 394
R1231 VSS.n2103 VSS.n250 394
R1232 VSS.n2103 VSS.n252 394
R1233 VSS.n2099 VSS.n252 394
R1234 VSS.n2099 VSS.n257 394
R1235 VSS.n2095 VSS.n257 394
R1236 VSS.n2095 VSS.n259 394
R1237 VSS.n2091 VSS.n259 394
R1238 VSS.n2091 VSS.n264 394
R1239 VSS.n2087 VSS.n264 394
R1240 VSS.n2087 VSS.n266 394
R1241 VSS.n2083 VSS.n266 394
R1242 VSS.n2083 VSS.n271 394
R1243 VSS.n2079 VSS.n271 394
R1244 VSS.n2079 VSS.n273 394
R1245 VSS.n2075 VSS.n273 394
R1246 VSS.n2075 VSS.n279 394
R1247 VSS.n2071 VSS.n279 394
R1248 VSS.n2071 VSS.n281 394
R1249 VSS.n2067 VSS.n281 394
R1250 VSS.n2067 VSS.n286 394
R1251 VSS.n2063 VSS.n286 394
R1252 VSS.n2063 VSS.n288 394
R1253 VSS.n2059 VSS.n288 394
R1254 VSS.n2059 VSS.n293 394
R1255 VSS.n2055 VSS.n293 394
R1256 VSS.n2055 VSS.n295 394
R1257 VSS.n2051 VSS.n295 394
R1258 VSS.n2051 VSS.n300 394
R1259 VSS.n2047 VSS.n300 394
R1260 VSS.n2047 VSS.n302 394
R1261 VSS.n2043 VSS.n302 394
R1262 VSS.n2043 VSS.n307 394
R1263 VSS.n2039 VSS.n307 394
R1264 VSS.n2039 VSS.n309 394
R1265 VSS.n2035 VSS.n309 394
R1266 VSS.n2035 VSS.n314 394
R1267 VSS.n2031 VSS.n314 394
R1268 VSS.n2031 VSS.n316 394
R1269 VSS.n2027 VSS.n316 394
R1270 VSS.n2027 VSS.n321 394
R1271 VSS.n2023 VSS.n321 394
R1272 VSS.n2023 VSS.n323 394
R1273 VSS.n2019 VSS.n323 394
R1274 VSS.n2019 VSS.n328 394
R1275 VSS.n2015 VSS.n328 394
R1276 VSS.n2015 VSS.n330 394
R1277 VSS.n2011 VSS.n330 394
R1278 VSS.n2011 VSS.n335 394
R1279 VSS.n2007 VSS.n335 394
R1280 VSS.n2007 VSS.n337 394
R1281 VSS.n2003 VSS.n337 394
R1282 VSS.n1829 VSS.n398 394
R1283 VSS.n1825 VSS.n1824 394
R1284 VSS.n1821 VSS.n1820 394
R1285 VSS.n1817 VSS.n1816 394
R1286 VSS.n1813 VSS.n1812 394
R1287 VSS.n1809 VSS.n1808 394
R1288 VSS.n1805 VSS.n1804 394
R1289 VSS.n1801 VSS.n1800 394
R1290 VSS.n1793 VSS.n1792 394
R1291 VSS.n1790 VSS.n1789 394
R1292 VSS.n406 VSS.n405 394
R1293 VSS.n1782 VSS.n1781 394
R1294 VSS.n1778 VSS.n1777 394
R1295 VSS.n1774 VSS.n1773 394
R1296 VSS.n1770 VSS.n1769 394
R1297 VSS.n1766 VSS.n1765 394
R1298 VSS.n1762 VSS.n1761 394
R1299 VSS.n1758 VSS.n1757 394
R1300 VSS.n1754 VSS.n379 394
R1301 VSS.n1837 VSS.n377 394
R1302 VSS.n1837 VSS.n372 394
R1303 VSS.n1846 VSS.n372 394
R1304 VSS.n1847 VSS.n1846 394
R1305 VSS.n1847 VSS.n240 394
R1306 VSS.n1850 VSS.n240 394
R1307 VSS.n1850 VSS.n247 394
R1308 VSS.n248 VSS.n247 394
R1309 VSS.n249 VSS.n248 394
R1310 VSS.n1855 VSS.n249 394
R1311 VSS.n1855 VSS.n254 394
R1312 VSS.n255 VSS.n254 394
R1313 VSS.n256 VSS.n255 394
R1314 VSS.n1860 VSS.n256 394
R1315 VSS.n1860 VSS.n261 394
R1316 VSS.n262 VSS.n261 394
R1317 VSS.n263 VSS.n262 394
R1318 VSS.n1865 VSS.n263 394
R1319 VSS.n1865 VSS.n268 394
R1320 VSS.n269 VSS.n268 394
R1321 VSS.n270 VSS.n269 394
R1322 VSS.n1870 VSS.n270 394
R1323 VSS.n1870 VSS.n275 394
R1324 VSS.n276 VSS.n275 394
R1325 VSS.n277 VSS.n276 394
R1326 VSS.n1875 VSS.n277 394
R1327 VSS.n1875 VSS.n282 394
R1328 VSS.n283 VSS.n282 394
R1329 VSS.n284 VSS.n283 394
R1330 VSS.n1880 VSS.n284 394
R1331 VSS.n1880 VSS.n289 394
R1332 VSS.n290 VSS.n289 394
R1333 VSS.n291 VSS.n290 394
R1334 VSS.n1885 VSS.n291 394
R1335 VSS.n1885 VSS.n296 394
R1336 VSS.n297 VSS.n296 394
R1337 VSS.n298 VSS.n297 394
R1338 VSS.n1890 VSS.n298 394
R1339 VSS.n1890 VSS.n303 394
R1340 VSS.n304 VSS.n303 394
R1341 VSS.n305 VSS.n304 394
R1342 VSS.n1895 VSS.n305 394
R1343 VSS.n1895 VSS.n310 394
R1344 VSS.n311 VSS.n310 394
R1345 VSS.n312 VSS.n311 394
R1346 VSS.n1900 VSS.n312 394
R1347 VSS.n1900 VSS.n317 394
R1348 VSS.n318 VSS.n317 394
R1349 VSS.n319 VSS.n318 394
R1350 VSS.n1905 VSS.n319 394
R1351 VSS.n1905 VSS.n324 394
R1352 VSS.n325 VSS.n324 394
R1353 VSS.n326 VSS.n325 394
R1354 VSS.n1910 VSS.n326 394
R1355 VSS.n1910 VSS.n331 394
R1356 VSS.n332 VSS.n331 394
R1357 VSS.n333 VSS.n332 394
R1358 VSS.n1915 VSS.n333 394
R1359 VSS.n1915 VSS.n338 394
R1360 VSS.n339 VSS.n338 394
R1361 VSS.n340 VSS.n339 394
R1362 VSS.n1999 VSS.n1997 394
R1363 VSS.n1997 VSS.n1996 394
R1364 VSS.n1993 VSS.n1992 394
R1365 VSS.n1990 VSS.n346 394
R1366 VSS.n1986 VSS.n1984 394
R1367 VSS.n1982 VSS.n348 394
R1368 VSS.n1978 VSS.n1976 394
R1369 VSS.n1974 VSS.n350 394
R1370 VSS.n1968 VSS.n1966 394
R1371 VSS.n1963 VSS.n1962 394
R1372 VSS.n1953 VSS.n1952 394
R1373 VSS.n1955 VSS.n1951 394
R1374 VSS.n1948 VSS.n1947 394
R1375 VSS.n1945 VSS.n365 394
R1376 VSS.n1941 VSS.n1939 394
R1377 VSS.n1937 VSS.n367 394
R1378 VSS.n1933 VSS.n1931 394
R1379 VSS.n1929 VSS.n369 394
R1380 VSS.n1925 VSS.n1923 394
R1381 VSS.n636 VSS.n55 394
R1382 VSS.n2558 VSS.n55 394
R1383 VSS.n2558 VSS.n53 394
R1384 VSS.n2562 VSS.n53 394
R1385 VSS.n2562 VSS.n48 394
R1386 VSS.n2570 VSS.n48 394
R1387 VSS.n2570 VSS.n46 394
R1388 VSS.n2574 VSS.n46 394
R1389 VSS.n2574 VSS.n39 394
R1390 VSS.n2600 VSS.n39 394
R1391 VSS.n2600 VSS.n37 394
R1392 VSS.n1540 VSS.n637 394
R1393 VSS.n1536 VSS.n1535 394
R1394 VSS.n1532 VSS.n1531 394
R1395 VSS.n1528 VSS.n1527 394
R1396 VSS.n1524 VSS.n1523 394
R1397 VSS.n1520 VSS.n1519 394
R1398 VSS.n1516 VSS.n1515 394
R1399 VSS.n1512 VSS.n1511 394
R1400 VSS.n1508 VSS.n1507 394
R1401 VSS.n1504 VSS.n1503 394
R1402 VSS.n1500 VSS.n1499 394
R1403 VSS.n1495 VSS.n642 394
R1404 VSS.n642 VSS.n56 394
R1405 VSS.n56 VSS.n51 394
R1406 VSS.n2564 VSS.n51 394
R1407 VSS.n2564 VSS.n49 394
R1408 VSS.n2568 VSS.n49 394
R1409 VSS.n2568 VSS.n43 394
R1410 VSS.n2576 VSS.n43 394
R1411 VSS.n2576 VSS.n40 394
R1412 VSS.n2598 VSS.n40 394
R1413 VSS.n2598 VSS.n41 394
R1414 VSS.n36 VSS.n35 394
R1415 VSS.n2617 VSS.n35 394
R1416 VSS.n2615 VSS.n2614 394
R1417 VSS.n2611 VSS.n2610 394
R1418 VSS.n2606 VSS.n2605 394
R1419 VSS.n29 VSS.n27 394
R1420 VSS.n2626 VSS.n19 394
R1421 VSS.n2580 VSS.n20 394
R1422 VSS.n2584 VSS.n2583 394
R1423 VSS.n2588 VSS.n2587 394
R1424 VSS.n2592 VSS.n2591 394
R1425 VSS.n1627 VSS.n573 394
R1426 VSS.n1623 VSS.n573 394
R1427 VSS.n1623 VSS.n576 394
R1428 VSS.n588 VSS.n576 394
R1429 VSS.n1613 VSS.n588 394
R1430 VSS.n1613 VSS.n589 394
R1431 VSS.n1609 VSS.n589 394
R1432 VSS.n1609 VSS.n592 394
R1433 VSS.n603 VSS.n592 394
R1434 VSS.n1599 VSS.n603 394
R1435 VSS.n1599 VSS.n604 394
R1436 VSS.n946 VSS.n572 394
R1437 VSS.n950 VSS.n948 394
R1438 VSS.n954 VSS.n943 394
R1439 VSS.n958 VSS.n956 394
R1440 VSS.n962 VSS.n941 394
R1441 VSS.n966 VSS.n964 394
R1442 VSS.n970 VSS.n939 394
R1443 VSS.n974 VSS.n972 394
R1444 VSS.n978 VSS.n937 394
R1445 VSS.n981 VSS.n980 394
R1446 VSS.n985 VSS.n984 394
R1447 VSS.n1067 VSS.n570 394
R1448 VSS.n1067 VSS.n577 394
R1449 VSS.n1061 VSS.n577 394
R1450 VSS.n1061 VSS.n1060 394
R1451 VSS.n1060 VSS.n587 394
R1452 VSS.n994 VSS.n587 394
R1453 VSS.n994 VSS.n594 394
R1454 VSS.n1051 VSS.n594 394
R1455 VSS.n1051 VSS.n1050 394
R1456 VSS.n1050 VSS.n601 394
R1457 VSS.n1551 VSS.n601 394
R1458 VSS.n1592 VSS.n607 394
R1459 VSS.n1592 VSS.n619 394
R1460 VSS.n1588 VSS.n1587 394
R1461 VSS.n1584 VSS.n1583 394
R1462 VSS.n1580 VSS.n1579 394
R1463 VSS.n1576 VSS.n1575 394
R1464 VSS.n1572 VSS.n1571 394
R1465 VSS.n1568 VSS.n1567 394
R1466 VSS.n1564 VSS.n1563 394
R1467 VSS.n1560 VSS.n1559 394
R1468 VSS.n1556 VSS.n1555 394
R1469 VSS.n1343 VSS.n716 394
R1470 VSS.n1358 VSS.n716 394
R1471 VSS.n1358 VSS.n714 394
R1472 VSS.n1362 VSS.n714 394
R1473 VSS.n1362 VSS.n703 394
R1474 VSS.n1417 VSS.n703 394
R1475 VSS.n1417 VSS.n704 394
R1476 VSS.n1413 VSS.n704 394
R1477 VSS.n1413 VSS.n707 394
R1478 VSS.n707 VSS.n508 394
R1479 VSS.n1643 VSS.n508 394
R1480 VSS.n1339 VSS.n1279 394
R1481 VSS.n1337 VSS.n1336 394
R1482 VSS.n1334 VSS.n1282 394
R1483 VSS.n1330 VSS.n1329 394
R1484 VSS.n1327 VSS.n1285 394
R1485 VSS.n1323 VSS.n1322 394
R1486 VSS.n1320 VSS.n1288 394
R1487 VSS.n1316 VSS.n1315 394
R1488 VSS.n1313 VSS.n1291 394
R1489 VSS.n1309 VSS.n1308 394
R1490 VSS.n1306 VSS.n1294 394
R1491 VSS.n1298 VSS.n1276 394
R1492 VSS.n1298 VSS.n717 394
R1493 VSS.n1295 VSS.n717 394
R1494 VSS.n1295 VSS.n712 394
R1495 VSS.n1366 VSS.n712 394
R1496 VSS.n1366 VSS.n701 394
R1497 VSS.n902 VSS.n701 394
R1498 VSS.n902 VSS.n709 394
R1499 VSS.n1375 VSS.n709 394
R1500 VSS.n1375 VSS.n505 394
R1501 VSS.n1645 VSS.n505 394
R1502 VSS.n1639 VSS.n512 394
R1503 VSS.n524 VSS.n512 394
R1504 VSS.n528 VSS.n527 394
R1505 VSS.n532 VSS.n531 394
R1506 VSS.n536 VSS.n535 394
R1507 VSS.n540 VSS.n539 394
R1508 VSS.n544 VSS.n543 394
R1509 VSS.n548 VSS.n547 394
R1510 VSS.n552 VSS.n551 394
R1511 VSS.n556 VSS.n555 394
R1512 VSS.n561 VSS.n523 394
R1513 VSS.n2141 VSS.n2134 394
R1514 VSS.n2139 VSS.n2138 394
R1515 VSS.n2145 VSS.n2128 394
R1516 VSS.n2153 VSS.n2128 394
R1517 VSS.n2153 VSS.n2126 394
R1518 VSS.n2157 VSS.n2126 394
R1519 VSS.n2157 VSS.n2120 394
R1520 VSS.n2166 VSS.n2120 394
R1521 VSS.n2166 VSS.n2118 394
R1522 VSS.n2170 VSS.n2118 394
R1523 VSS.n2170 VSS.n234 394
R1524 VSS.n2178 VSS.n234 394
R1525 VSS.n2178 VSS.n232 394
R1526 VSS.n2182 VSS.n232 394
R1527 VSS.n2182 VSS.n226 394
R1528 VSS.n2190 VSS.n226 394
R1529 VSS.n2190 VSS.n224 394
R1530 VSS.n2194 VSS.n224 394
R1531 VSS.n2194 VSS.n218 394
R1532 VSS.n2202 VSS.n218 394
R1533 VSS.n2202 VSS.n216 394
R1534 VSS.n2206 VSS.n216 394
R1535 VSS.n2206 VSS.n210 394
R1536 VSS.n2214 VSS.n210 394
R1537 VSS.n2214 VSS.n208 394
R1538 VSS.n2218 VSS.n208 394
R1539 VSS.n2218 VSS.n202 394
R1540 VSS.n2226 VSS.n202 394
R1541 VSS.n2226 VSS.n200 394
R1542 VSS.n2230 VSS.n200 394
R1543 VSS.n2230 VSS.n193 394
R1544 VSS.n2238 VSS.n193 394
R1545 VSS.n2238 VSS.n191 394
R1546 VSS.n2242 VSS.n191 394
R1547 VSS.n2242 VSS.n185 394
R1548 VSS.n2250 VSS.n185 394
R1549 VSS.n2250 VSS.n183 394
R1550 VSS.n2254 VSS.n183 394
R1551 VSS.n2254 VSS.n177 394
R1552 VSS.n2262 VSS.n177 394
R1553 VSS.n2262 VSS.n175 394
R1554 VSS.n2266 VSS.n175 394
R1555 VSS.n2266 VSS.n169 394
R1556 VSS.n2274 VSS.n169 394
R1557 VSS.n2274 VSS.n167 394
R1558 VSS.n2278 VSS.n167 394
R1559 VSS.n2278 VSS.n161 394
R1560 VSS.n2286 VSS.n161 394
R1561 VSS.n2286 VSS.n159 394
R1562 VSS.n2290 VSS.n159 394
R1563 VSS.n2290 VSS.n153 394
R1564 VSS.n2299 VSS.n153 394
R1565 VSS.n2299 VSS.n151 394
R1566 VSS.n2303 VSS.n151 394
R1567 VSS.n2303 VSS.n140 394
R1568 VSS.n2311 VSS.n141 394
R1569 VSS.n2311 VSS.n145 394
R1570 VSS.n2147 VSS.n2130 394
R1571 VSS.n2151 VSS.n2130 394
R1572 VSS.n2151 VSS.n2124 394
R1573 VSS.n2159 VSS.n2124 394
R1574 VSS.n2159 VSS.n2122 394
R1575 VSS.n2163 VSS.n2122 394
R1576 VSS.n2163 VSS.n238 394
R1577 VSS.n2172 VSS.n238 394
R1578 VSS.n2172 VSS.n236 394
R1579 VSS.n2176 VSS.n236 394
R1580 VSS.n2176 VSS.n230 394
R1581 VSS.n2184 VSS.n230 394
R1582 VSS.n2184 VSS.n228 394
R1583 VSS.n2188 VSS.n228 394
R1584 VSS.n2188 VSS.n222 394
R1585 VSS.n2196 VSS.n222 394
R1586 VSS.n2196 VSS.n220 394
R1587 VSS.n2200 VSS.n220 394
R1588 VSS.n2200 VSS.n214 394
R1589 VSS.n2208 VSS.n214 394
R1590 VSS.n2208 VSS.n212 394
R1591 VSS.n2212 VSS.n212 394
R1592 VSS.n2212 VSS.n206 394
R1593 VSS.n2220 VSS.n206 394
R1594 VSS.n2220 VSS.n204 394
R1595 VSS.n2224 VSS.n204 394
R1596 VSS.n2224 VSS.n197 394
R1597 VSS.n2232 VSS.n197 394
R1598 VSS.n2232 VSS.n195 394
R1599 VSS.n2236 VSS.n195 394
R1600 VSS.n2236 VSS.n189 394
R1601 VSS.n2244 VSS.n189 394
R1602 VSS.n2244 VSS.n187 394
R1603 VSS.n2248 VSS.n187 394
R1604 VSS.n2248 VSS.n181 394
R1605 VSS.n2256 VSS.n181 394
R1606 VSS.n2256 VSS.n179 394
R1607 VSS.n2260 VSS.n179 394
R1608 VSS.n2260 VSS.n173 394
R1609 VSS.n2268 VSS.n173 394
R1610 VSS.n2268 VSS.n171 394
R1611 VSS.n2272 VSS.n171 394
R1612 VSS.n2272 VSS.n165 394
R1613 VSS.n2280 VSS.n165 394
R1614 VSS.n2280 VSS.n163 394
R1615 VSS.n2284 VSS.n163 394
R1616 VSS.n2284 VSS.n157 394
R1617 VSS.n2292 VSS.n157 394
R1618 VSS.n2292 VSS.n155 394
R1619 VSS.n2297 VSS.n155 394
R1620 VSS.n2297 VSS.n148 394
R1621 VSS.n2305 VSS.n148 394
R1622 VSS.n2306 VSS.n2305 394
R1623 VSS.n1091 VSS.n771 394
R1624 VSS.n1087 VSS.n771 394
R1625 VSS.n1087 VSS.n773 394
R1626 VSS.n900 VSS.n773 394
R1627 VSS.n905 VSS.n900 394
R1628 VSS.n905 VSS.n897 394
R1629 VSS.n911 VSS.n897 394
R1630 VSS.n911 VSS.n895 394
R1631 VSS.n915 VSS.n895 394
R1632 VSS.n917 VSS.n915 394
R1633 VSS.n917 VSS.n893 394
R1634 VSS.n921 VSS.n893 394
R1635 VSS.n921 VSS.n891 394
R1636 VSS.n925 VSS.n891 394
R1637 VSS.n925 VSS.n888 394
R1638 VSS.n932 VSS.n888 394
R1639 VSS.n932 VSS.n889 394
R1640 VSS.n889 VSS.n884 394
R1641 VSS.n1074 VSS.n884 394
R1642 VSS.n1074 VSS.n885 394
R1643 VSS.n1017 VSS.n885 394
R1644 VSS.n1023 VSS.n1017 394
R1645 VSS.n1023 VSS.n1019 394
R1646 VSS.n1019 VSS.n1004 394
R1647 VSS.n1047 VSS.n1004 394
R1648 VSS.n1047 VSS.n1005 394
R1649 VSS.n1043 VSS.n1005 394
R1650 VSS.n1043 VSS.n1040 394
R1651 VSS.n1040 VSS.n1039 394
R1652 VSS.n1039 VSS.n1008 394
R1653 VSS.n1035 VSS.n1008 394
R1654 VSS.n1035 VSS.n1011 394
R1655 VSS.n1011 VSS.n124 394
R1656 VSS.n2352 VSS.n124 394
R1657 VSS.n2352 VSS.n120 394
R1658 VSS.n2356 VSS.n120 394
R1659 VSS.n2356 VSS.n122 394
R1660 VSS.n122 VSS.n116 394
R1661 VSS.n115 VSS.n114 394
R1662 VSS.n2391 VSS.n114 394
R1663 VSS.n2389 VSS.n2388 394
R1664 VSS.n2385 VSS.n2384 394
R1665 VSS.n2381 VSS.n2380 394
R1666 VSS.n2377 VSS.n2376 394
R1667 VSS.n2373 VSS.n2372 394
R1668 VSS.n2369 VSS.n2368 394
R1669 VSS.n2365 VSS.n2364 394
R1670 VSS.n2399 VSS.n103 394
R1671 VSS.n2400 VSS.n2399 394
R1672 VSS.n2402 VSS.n101 394
R1673 VSS.n2410 VSS.n2408 394
R1674 VSS.n2414 VSS.n99 394
R1675 VSS.n2418 VSS.n2416 394
R1676 VSS.n2422 VSS.n97 394
R1677 VSS.n2426 VSS.n2424 394
R1678 VSS.n2430 VSS.n95 394
R1679 VSS.n2434 VSS.n2432 394
R1680 VSS.n2438 VSS.n93 394
R1681 VSS.n2442 VSS.n2440 394
R1682 VSS.n2446 VSS.n91 394
R1683 VSS.n2450 VSS.n2448 394
R1684 VSS.n2458 VSS.n2456 394
R1685 VSS.n2462 VSS.n87 394
R1686 VSS.n2466 VSS.n2464 394
R1687 VSS.n2470 VSS.n85 394
R1688 VSS.n2474 VSS.n2472 394
R1689 VSS.n2478 VSS.n83 394
R1690 VSS.n2482 VSS.n2480 394
R1691 VSS.n2486 VSS.n81 394
R1692 VSS.n2490 VSS.n2488 394
R1693 VSS.n2494 VSS.n79 394
R1694 VSS.n2498 VSS.n2496 394
R1695 VSS.n2506 VSS.n2504 394
R1696 VSS.n2510 VSS.n75 394
R1697 VSS.n2514 VSS.n2512 394
R1698 VSS.n2518 VSS.n73 394
R1699 VSS.n2522 VSS.n2520 394
R1700 VSS.n2526 VSS.n71 394
R1701 VSS.n2530 VSS.n2528 394
R1702 VSS.n2534 VSS.n69 394
R1703 VSS.n2538 VSS.n2536 394
R1704 VSS.n2542 VSS.n67 394
R1705 VSS.n2545 VSS.n2544 394
R1706 VSS.n1355 VSS.n719 394
R1707 VSS.n1355 VSS.n720 394
R1708 VSS.n720 VSS.n699 394
R1709 VSS.n1420 VSS.n699 394
R1710 VSS.n1420 VSS.n700 394
R1711 VSS.n1377 VSS.n700 394
R1712 VSS.n1410 VSS.n1377 394
R1713 VSS.n1410 VSS.n1380 394
R1714 VSS.n1385 VSS.n1380 394
R1715 VSS.n1385 VSS.n1384 394
R1716 VSS.n1384 VSS.n564 394
R1717 VSS.n1635 VSS.n564 394
R1718 VSS.n1635 VSS.n565 394
R1719 VSS.n1631 VSS.n565 394
R1720 VSS.n1631 VSS.n568 394
R1721 VSS.n1397 VSS.n568 394
R1722 VSS.n1397 VSS.n579 394
R1723 VSS.n1620 VSS.n579 394
R1724 VSS.n1620 VSS.n580 394
R1725 VSS.n1616 VSS.n580 394
R1726 VSS.n1616 VSS.n584 394
R1727 VSS.n596 VSS.n584 394
R1728 VSS.n1606 VSS.n596 394
R1729 VSS.n1606 VSS.n597 394
R1730 VSS.n1602 VSS.n597 394
R1731 VSS.n1602 VSS.n600 394
R1732 VSS.n1548 VSS.n600 394
R1733 VSS.n1548 VSS.n621 394
R1734 VSS.n1544 VSS.n621 394
R1735 VSS.n1544 VSS.n623 394
R1736 VSS.n648 VSS.n623 394
R1737 VSS.n648 VSS.n646 394
R1738 VSS.n1492 VSS.n646 394
R1739 VSS.n1492 VSS.n58 394
R1740 VSS.n2555 VSS.n58 394
R1741 VSS.n2555 VSS.n60 394
R1742 VSS.n65 VSS.n60 394
R1743 VSS.n2548 VSS.n65 394
R1744 VSS.n1097 VSS.n769 394
R1745 VSS.n1101 VSS.n1099 394
R1746 VSS.n1105 VSS.n767 394
R1747 VSS.n1109 VSS.n1107 394
R1748 VSS.n1113 VSS.n765 394
R1749 VSS.n1117 VSS.n1115 394
R1750 VSS.n1121 VSS.n763 394
R1751 VSS.n1125 VSS.n1123 394
R1752 VSS.n1129 VSS.n761 394
R1753 VSS.n1132 VSS.n1131 394
R1754 VSS.n1136 VSS.n1135 394
R1755 VSS.n1140 VSS.n1139 394
R1756 VSS.n1144 VSS.n1143 394
R1757 VSS.n1148 VSS.n1147 394
R1758 VSS.n1152 VSS.n1151 394
R1759 VSS.n1156 VSS.n1155 394
R1760 VSS.n1160 VSS.n1159 394
R1761 VSS.n1164 VSS.n1163 394
R1762 VSS.n1168 VSS.n1167 394
R1763 VSS.n1172 VSS.n1171 394
R1764 VSS.n1176 VSS.n1175 394
R1765 VSS.n1180 VSS.n1179 394
R1766 VSS.n1184 VSS.n1183 394
R1767 VSS.n1188 VSS.n1187 394
R1768 VSS.n1192 VSS.n1191 394
R1769 VSS.n1196 VSS.n1195 394
R1770 VSS.n1200 VSS.n1199 394
R1771 VSS.n1204 VSS.n1203 394
R1772 VSS.n1208 VSS.n1207 394
R1773 VSS.n1212 VSS.n1211 394
R1774 VSS.n1216 VSS.n1215 394
R1775 VSS.n1220 VSS.n1219 394
R1776 VSS.n1224 VSS.n1223 394
R1777 VSS.n1228 VSS.n1227 394
R1778 VSS.n1232 VSS.n1231 394
R1779 VSS.n1236 VSS.n1235 394
R1780 VSS.n1240 VSS.n1239 394
R1781 VSS.n1244 VSS.n1243 394
R1782 VSS.n1248 VSS.n1247 394
R1783 VSS.n1252 VSS.n1251 394
R1784 VSS.n1256 VSS.n1255 394
R1785 VSS.n1260 VSS.n1259 394
R1786 VSS.n1264 VSS.n1263 394
R1787 VSS.n1268 VSS.n1267 394
R1788 VSS.n1270 VSS.n759 394
R1789 VSS.n1274 VSS.n722 394
R1790 VSS.n2231 VSS.n194 328.791
R1791 VSS.n2237 VSS.n194 328.791
R1792 VSS.n2237 VSS.n190 328.791
R1793 VSS.n2243 VSS.n190 328.791
R1794 VSS.n2243 VSS.n186 328.791
R1795 VSS.n2249 VSS.n186 328.791
R1796 VSS.n2249 VSS.n182 328.791
R1797 VSS.n2255 VSS.n182 328.791
R1798 VSS.n2255 VSS.n178 328.791
R1799 VSS.n2261 VSS.n178 328.791
R1800 VSS.n2261 VSS.n174 328.791
R1801 VSS.n2267 VSS.n174 328.791
R1802 VSS.n2267 VSS.n170 328.791
R1803 VSS.n2273 VSS.n170 328.791
R1804 VSS.n2273 VSS.n166 328.791
R1805 VSS.n2279 VSS.n166 328.791
R1806 VSS.n2279 VSS.n162 328.791
R1807 VSS.n2285 VSS.n162 328.791
R1808 VSS.n2285 VSS.n158 328.791
R1809 VSS.n2291 VSS.n158 328.791
R1810 VSS.n2291 VSS.n154 328.791
R1811 VSS.n2298 VSS.n154 328.791
R1812 VSS.n2298 VSS.n150 328.791
R1813 VSS.n2304 VSS.n150 328.791
R1814 VSS.n2304 VSS.n142 328.791
R1815 VSS.n477 VSS.n476 325.69
R1816 VSS.n422 VSS.n417 325.69
R1817 VSS.n1136 VSS.n725 269.089
R1818 VSS.n1139 VSS.n725 269.089
R1819 VSS.n723 VSS.n341 261
R1820 VSS.n1481 VSS.t71 259.252
R1821 VSS.n1432 VSS.t74 259.252
R1822 VSS.n776 VSS.t67 259.252
R1823 VSS.n126 VSS.t109 259.252
R1824 VSS.n1428 VSS.t107 258.99
R1825 VSS.n1429 VSS.t131 258.99
R1826 VSS.n1430 VSS.t65 258.99
R1827 VSS.n1431 VSS.t69 258.99
R1828 VSS.n654 VSS.t119 258.99
R1829 VSS.n1424 VSS.t99 258.99
R1830 VSS.n1425 VSS.t101 258.99
R1831 VSS.n1426 VSS.t105 258.99
R1832 VSS.n791 VSS.t117 258.99
R1833 VSS.n790 VSS.t121 258.99
R1834 VSS.n789 VSS.t103 258.99
R1835 VSS.n788 VSS.t82 258.99
R1836 VSS.n784 VSS.t112 258.99
R1837 VSS.n785 VSS.t97 258.99
R1838 VSS.n786 VSS.t80 258.99
R1839 VSS.n787 VSS.t129 258.99
R1840 VSS.n689 VSS.n688 253.042
R1841 VSS.n1444 VSS.n1442 253.042
R1842 VSS.n825 VSS.n795 253.042
R1843 VSS.n852 VSS.n851 253.042
R1844 VSS.n2137 VSS.n2133 218.815
R1845 VSS.n2140 VSS.n2133 218.815
R1846 VSS.n2313 VSS.n2312 218.815
R1847 VSS.n2312 VSS.n143 218.815
R1848 VSS.n1638 VSS.n1637 218.815
R1849 VSS.n1637 VSS.n514 218.815
R1850 VSS.n1637 VSS.n515 218.815
R1851 VSS.n1637 VSS.n516 218.815
R1852 VSS.n1637 VSS.n517 218.815
R1853 VSS.n1637 VSS.n518 218.815
R1854 VSS.n1637 VSS.n519 218.815
R1855 VSS.n1637 VSS.n520 218.815
R1856 VSS.n1637 VSS.n521 218.815
R1857 VSS.n1637 VSS.n522 218.815
R1858 VSS.n1637 VSS.n562 218.815
R1859 VSS.n1301 VSS.n723 218.815
R1860 VSS.n1307 VSS.n723 218.815
R1861 VSS.n1293 VSS.n723 218.815
R1862 VSS.n1314 VSS.n723 218.815
R1863 VSS.n1290 VSS.n723 218.815
R1864 VSS.n1321 VSS.n723 218.815
R1865 VSS.n1287 VSS.n723 218.815
R1866 VSS.n1328 VSS.n723 218.815
R1867 VSS.n1284 VSS.n723 218.815
R1868 VSS.n1335 VSS.n723 218.815
R1869 VSS.n1338 VSS.n723 218.815
R1870 VSS.n1594 VSS.n1593 218.815
R1871 VSS.n1593 VSS.n609 218.815
R1872 VSS.n1593 VSS.n610 218.815
R1873 VSS.n1593 VSS.n611 218.815
R1874 VSS.n1593 VSS.n612 218.815
R1875 VSS.n1593 VSS.n613 218.815
R1876 VSS.n1593 VSS.n614 218.815
R1877 VSS.n1593 VSS.n615 218.815
R1878 VSS.n1593 VSS.n616 218.815
R1879 VSS.n1593 VSS.n617 218.815
R1880 VSS.n1593 VSS.n618 218.815
R1881 VSS.n986 VSS.n569 218.815
R1882 VSS.n935 VSS.n569 218.815
R1883 VSS.n979 VSS.n569 218.815
R1884 VSS.n973 VSS.n569 218.815
R1885 VSS.n971 VSS.n569 218.815
R1886 VSS.n965 VSS.n569 218.815
R1887 VSS.n963 VSS.n569 218.815
R1888 VSS.n957 VSS.n569 218.815
R1889 VSS.n955 VSS.n569 218.815
R1890 VSS.n949 VSS.n569 218.815
R1891 VSS.n947 VSS.n569 218.815
R1892 VSS.n2624 VSS.n2623 218.815
R1893 VSS.n2624 VSS.n22 218.815
R1894 VSS.n2624 VSS.n23 218.815
R1895 VSS.n2624 VSS.n24 218.815
R1896 VSS.n2624 VSS.n25 218.815
R1897 VSS.n2624 VSS.n30 218.815
R1898 VSS.n2625 VSS.n2624 218.815
R1899 VSS.n2624 VSS.n31 218.815
R1900 VSS.n2624 VSS.n32 218.815
R1901 VSS.n2624 VSS.n33 218.815
R1902 VSS.n2624 VSS.n34 218.815
R1903 VSS.n1541 VSS.n625 218.815
R1904 VSS.n1541 VSS.n626 218.815
R1905 VSS.n1541 VSS.n627 218.815
R1906 VSS.n1541 VSS.n628 218.815
R1907 VSS.n1541 VSS.n629 218.815
R1908 VSS.n1541 VSS.n630 218.815
R1909 VSS.n1541 VSS.n631 218.815
R1910 VSS.n1541 VSS.n632 218.815
R1911 VSS.n1541 VSS.n633 218.815
R1912 VSS.n1541 VSS.n634 218.815
R1913 VSS.n1541 VSS.n635 218.815
R1914 VSS.n1998 VSS.n341 218.815
R1915 VSS.n344 VSS.n341 218.815
R1916 VSS.n1991 VSS.n341 218.815
R1917 VSS.n1985 VSS.n341 218.815
R1918 VSS.n1983 VSS.n341 218.815
R1919 VSS.n1977 VSS.n341 218.815
R1920 VSS.n1975 VSS.n341 218.815
R1921 VSS.n1967 VSS.n341 218.815
R1922 VSS.n354 VSS.n341 218.815
R1923 VSS.n356 VSS.n341 218.815
R1924 VSS.n1954 VSS.n341 218.815
R1925 VSS.n362 VSS.n341 218.815
R1926 VSS.n1946 VSS.n341 218.815
R1927 VSS.n1940 VSS.n341 218.815
R1928 VSS.n1938 VSS.n341 218.815
R1929 VSS.n1932 VSS.n341 218.815
R1930 VSS.n1930 VSS.n341 218.815
R1931 VSS.n1924 VSS.n341 218.815
R1932 VSS.n1922 VSS.n341 218.815
R1933 VSS.n1831 VSS.n1830 218.815
R1934 VSS.n1830 VSS.n380 218.815
R1935 VSS.n1830 VSS.n381 218.815
R1936 VSS.n1830 VSS.n382 218.815
R1937 VSS.n1830 VSS.n383 218.815
R1938 VSS.n1830 VSS.n384 218.815
R1939 VSS.n1830 VSS.n385 218.815
R1940 VSS.n1830 VSS.n386 218.815
R1941 VSS.n1830 VSS.n387 218.815
R1942 VSS.n1830 VSS.n388 218.815
R1943 VSS.n1830 VSS.n389 218.815
R1944 VSS.n1830 VSS.n390 218.815
R1945 VSS.n1830 VSS.n391 218.815
R1946 VSS.n1830 VSS.n392 218.815
R1947 VSS.n1830 VSS.n393 218.815
R1948 VSS.n1830 VSS.n394 218.815
R1949 VSS.n1830 VSS.n395 218.815
R1950 VSS.n1830 VSS.n396 218.815
R1951 VSS.n1830 VSS.n397 218.815
R1952 VSS.n1346 VSS.n1345 218.815
R1953 VSS.n1345 VSS.n1275 218.815
R1954 VSS.n1345 VSS.n758 218.815
R1955 VSS.n1345 VSS.n757 218.815
R1956 VSS.n1345 VSS.n756 218.815
R1957 VSS.n1345 VSS.n755 218.815
R1958 VSS.n1345 VSS.n754 218.815
R1959 VSS.n1345 VSS.n753 218.815
R1960 VSS.n1345 VSS.n752 218.815
R1961 VSS.n1345 VSS.n751 218.815
R1962 VSS.n1345 VSS.n750 218.815
R1963 VSS.n1345 VSS.n748 218.815
R1964 VSS.n1345 VSS.n747 218.815
R1965 VSS.n1345 VSS.n746 218.815
R1966 VSS.n1345 VSS.n745 218.815
R1967 VSS.n1345 VSS.n744 218.815
R1968 VSS.n1345 VSS.n743 218.815
R1969 VSS.n1345 VSS.n742 218.815
R1970 VSS.n1345 VSS.n741 218.815
R1971 VSS.n1345 VSS.n740 218.815
R1972 VSS.n1345 VSS.n739 218.815
R1973 VSS.n1345 VSS.n738 218.815
R1974 VSS.n1345 VSS.n736 218.815
R1975 VSS.n1345 VSS.n735 218.815
R1976 VSS.n1345 VSS.n734 218.815
R1977 VSS.n1345 VSS.n733 218.815
R1978 VSS.n1345 VSS.n732 218.815
R1979 VSS.n1345 VSS.n731 218.815
R1980 VSS.n1345 VSS.n730 218.815
R1981 VSS.n1345 VSS.n729 218.815
R1982 VSS.n1345 VSS.n728 218.815
R1983 VSS.n1345 VSS.n727 218.815
R1984 VSS.n1345 VSS.n726 218.815
R1985 VSS.n1345 VSS.n724 218.815
R1986 VSS.n1130 VSS.n144 218.815
R1987 VSS.n1124 VSS.n144 218.815
R1988 VSS.n1122 VSS.n144 218.815
R1989 VSS.n1116 VSS.n144 218.815
R1990 VSS.n1114 VSS.n144 218.815
R1991 VSS.n1108 VSS.n144 218.815
R1992 VSS.n1106 VSS.n144 218.815
R1993 VSS.n1100 VSS.n144 218.815
R1994 VSS.n1098 VSS.n144 218.815
R1995 VSS.n1092 VSS.n144 218.815
R1996 VSS.n2398 VSS.n2397 218.815
R1997 VSS.n2398 VSS.n106 218.815
R1998 VSS.n2398 VSS.n107 218.815
R1999 VSS.n2398 VSS.n108 218.815
R2000 VSS.n2398 VSS.n109 218.815
R2001 VSS.n2398 VSS.n110 218.815
R2002 VSS.n2398 VSS.n111 218.815
R2003 VSS.n2398 VSS.n112 218.815
R2004 VSS.n2398 VSS.n113 218.815
R2005 VSS.n2401 VSS.n44 218.815
R2006 VSS.n2407 VSS.n44 218.815
R2007 VSS.n2409 VSS.n44 218.815
R2008 VSS.n2415 VSS.n44 218.815
R2009 VSS.n2417 VSS.n44 218.815
R2010 VSS.n2423 VSS.n44 218.815
R2011 VSS.n2425 VSS.n44 218.815
R2012 VSS.n2431 VSS.n44 218.815
R2013 VSS.n2433 VSS.n44 218.815
R2014 VSS.n2439 VSS.n44 218.815
R2015 VSS.n2441 VSS.n44 218.815
R2016 VSS.n2447 VSS.n44 218.815
R2017 VSS.n2449 VSS.n44 218.815
R2018 VSS.n2455 VSS.n44 218.815
R2019 VSS.n2457 VSS.n44 218.815
R2020 VSS.n2463 VSS.n44 218.815
R2021 VSS.n2465 VSS.n44 218.815
R2022 VSS.n2471 VSS.n44 218.815
R2023 VSS.n2473 VSS.n44 218.815
R2024 VSS.n2479 VSS.n44 218.815
R2025 VSS.n2481 VSS.n44 218.815
R2026 VSS.n2487 VSS.n44 218.815
R2027 VSS.n2489 VSS.n44 218.815
R2028 VSS.n2495 VSS.n44 218.815
R2029 VSS.n2497 VSS.n44 218.815
R2030 VSS.n2503 VSS.n44 218.815
R2031 VSS.n2505 VSS.n44 218.815
R2032 VSS.n2511 VSS.n44 218.815
R2033 VSS.n2513 VSS.n44 218.815
R2034 VSS.n2519 VSS.n44 218.815
R2035 VSS.n2521 VSS.n44 218.815
R2036 VSS.n2527 VSS.n44 218.815
R2037 VSS.n2529 VSS.n44 218.815
R2038 VSS.n2535 VSS.n44 218.815
R2039 VSS.n2537 VSS.n44 218.815
R2040 VSS.n2543 VSS.n44 218.815
R2041 VSS.n1184 VSS.n737 198.87
R2042 VSS.n1232 VSS.n749 198.87
R2043 VSS.n1235 VSS.n749 198.87
R2044 VSS.n1187 VSS.n737 198.87
R2045 VSS.n1345 VSS.n749 193.066
R2046 VSS.n1345 VSS.n737 193.066
R2047 VSS.n2146 VSS.n2133 185.895
R2048 VSS.n667 VSS.n666 185
R2049 VSS.n672 VSS.n671 185
R2050 VSS.n674 VSS.n673 185
R2051 VSS.n663 VSS.n662 185
R2052 VSS.n680 VSS.n679 185
R2053 VSS.n682 VSS.n681 185
R2054 VSS.n659 VSS.n658 185
R2055 VSS.n688 VSS.n687 185
R2056 VSS.n1466 VSS.n1465 185
R2057 VSS.n1435 VSS.n1434 185
R2058 VSS.n1460 VSS.n1459 185
R2059 VSS.n1458 VSS.n1457 185
R2060 VSS.n1439 VSS.n1438 185
R2061 VSS.n1452 VSS.n1451 185
R2062 VSS.n1450 VSS.n1449 185
R2063 VSS.n1443 VSS.n1442 185
R2064 VSS.n826 VSS.n825 185
R2065 VSS.n824 VSS.n823 185
R2066 VSS.n799 VSS.n798 185
R2067 VSS.n818 VSS.n817 185
R2068 VSS.n816 VSS.n815 185
R2069 VSS.n803 VSS.n802 185
R2070 VSS.n810 VSS.n809 185
R2071 VSS.n808 VSS.n807 185
R2072 VSS.n853 VSS.n852 185
R2073 VSS.n848 VSS.n847 185
R2074 VSS.n859 VSS.n858 185
R2075 VSS.n861 VSS.n860 185
R2076 VSS.n844 VSS.n843 185
R2077 VSS.n868 VSS.n867 185
R2078 VSS.n870 VSS.n869 185
R2079 VSS.n872 VSS.n840 185
R2080 VSS.n476 VSS.n475 185
R2081 VSS.n453 VSS.n452 185
R2082 VSS.n470 VSS.n469 185
R2083 VSS.n464 VSS.n463 185
R2084 VSS.n464 VSS.n456 185
R2085 VSS.n436 VSS.n435 185
R2086 VSS.n435 VSS.n434 185
R2087 VSS.n422 VSS.n421 185
R2088 VSS.n424 VSS.n423 185
R2089 VSS.n426 VSS.n414 185
R2090 VSS.n1687 VSS.n1686 185
R2091 VSS.n1687 VSS.n1659 185
R2092 VSS.n1689 VSS.n1688 185
R2093 VSS.n1688 VSS.n1657 185
R2094 VSS.n1671 VSS.n1663 185
R2095 VSS.n1671 VSS.n1662 185
R2096 VSS.n1672 VSS.n1671 185
R2097 VSS.n1749 VSS.n1748 185
R2098 VSS.n1748 VSS.n1732 185
R2099 VSS.n1747 VSS.n1746 185
R2100 VSS.n1747 VSS.n1734 185
R2101 VSS.n1726 VSS.n1718 185
R2102 VSS.n1726 VSS.n1717 185
R2103 VSS.n1727 VSS.n1726 185
R2104 VSS.n668 VSS.t73 178.418
R2105 VSS.t75 VSS.n1433 178.418
R2106 VSS.n806 VSS.t111 178.418
R2107 VSS.t68 VSS.n873 178.418
R2108 VSS.t116 VSS.n468 175.332
R2109 VSS.t126 VSS.n427 175.332
R2110 VSS.n1090 VSS.n144 163.94
R2111 VSS.n2398 VSS.n105 163.94
R2112 VSS.n1345 VSS.n725 157.957
R2113 VSS.n1825 VSS.n397 147.374
R2114 VSS.n1821 VSS.n396 147.374
R2115 VSS.n1817 VSS.n395 147.374
R2116 VSS.n1813 VSS.n394 147.374
R2117 VSS.n1809 VSS.n393 147.374
R2118 VSS.n1805 VSS.n392 147.374
R2119 VSS.n1801 VSS.n391 147.374
R2120 VSS.n1792 VSS.n390 147.374
R2121 VSS.n1790 VSS.n389 147.374
R2122 VSS.n405 VSS.n388 147.374
R2123 VSS.n1782 VSS.n387 147.374
R2124 VSS.n1778 VSS.n386 147.374
R2125 VSS.n1774 VSS.n385 147.374
R2126 VSS.n1770 VSS.n384 147.374
R2127 VSS.n1766 VSS.n383 147.374
R2128 VSS.n1762 VSS.n382 147.374
R2129 VSS.n1758 VSS.n381 147.374
R2130 VSS.n1754 VSS.n380 147.374
R2131 VSS.n1832 VSS.n1831 147.374
R2132 VSS.n1998 VSS.n342 147.374
R2133 VSS.n1996 VSS.n344 147.374
R2134 VSS.n1992 VSS.n1991 147.374
R2135 VSS.n1985 VSS.n346 147.374
R2136 VSS.n1984 VSS.n1983 147.374
R2137 VSS.n1977 VSS.n348 147.374
R2138 VSS.n1976 VSS.n1975 147.374
R2139 VSS.n1967 VSS.n350 147.374
R2140 VSS.n1966 VSS.n354 147.374
R2141 VSS.n1962 VSS.n356 147.374
R2142 VSS.n1954 VSS.n1953 147.374
R2143 VSS.n1951 VSS.n362 147.374
R2144 VSS.n1947 VSS.n1946 147.374
R2145 VSS.n1940 VSS.n365 147.374
R2146 VSS.n1939 VSS.n1938 147.374
R2147 VSS.n1932 VSS.n367 147.374
R2148 VSS.n1931 VSS.n1930 147.374
R2149 VSS.n1924 VSS.n369 147.374
R2150 VSS.n1923 VSS.n1922 147.374
R2151 VSS.n1536 VSS.n635 147.374
R2152 VSS.n1532 VSS.n634 147.374
R2153 VSS.n1528 VSS.n633 147.374
R2154 VSS.n1524 VSS.n632 147.374
R2155 VSS.n1520 VSS.n631 147.374
R2156 VSS.n1516 VSS.n630 147.374
R2157 VSS.n1512 VSS.n629 147.374
R2158 VSS.n1508 VSS.n628 147.374
R2159 VSS.n1504 VSS.n627 147.374
R2160 VSS.n1500 VSS.n626 147.374
R2161 VSS.n1496 VSS.n625 147.374
R2162 VSS.n2623 VSS.n2622 147.374
R2163 VSS.n2617 VSS.n22 147.374
R2164 VSS.n2614 VSS.n23 147.374
R2165 VSS.n2610 VSS.n24 147.374
R2166 VSS.n2605 VSS.n25 147.374
R2167 VSS.n30 VSS.n29 147.374
R2168 VSS.n2626 VSS.n2625 147.374
R2169 VSS.n2580 VSS.n31 147.374
R2170 VSS.n2584 VSS.n32 147.374
R2171 VSS.n2588 VSS.n33 147.374
R2172 VSS.n2592 VSS.n34 147.374
R2173 VSS.n948 VSS.n947 147.374
R2174 VSS.n949 VSS.n943 147.374
R2175 VSS.n956 VSS.n955 147.374
R2176 VSS.n957 VSS.n941 147.374
R2177 VSS.n964 VSS.n963 147.374
R2178 VSS.n965 VSS.n939 147.374
R2179 VSS.n972 VSS.n971 147.374
R2180 VSS.n973 VSS.n937 147.374
R2181 VSS.n980 VSS.n979 147.374
R2182 VSS.n984 VSS.n935 147.374
R2183 VSS.n987 VSS.n986 147.374
R2184 VSS.n1595 VSS.n1594 147.374
R2185 VSS.n619 VSS.n609 147.374
R2186 VSS.n1587 VSS.n610 147.374
R2187 VSS.n1583 VSS.n611 147.374
R2188 VSS.n1579 VSS.n612 147.374
R2189 VSS.n1575 VSS.n613 147.374
R2190 VSS.n1571 VSS.n614 147.374
R2191 VSS.n1567 VSS.n615 147.374
R2192 VSS.n1563 VSS.n616 147.374
R2193 VSS.n1559 VSS.n617 147.374
R2194 VSS.n1555 VSS.n618 147.374
R2195 VSS.n1338 VSS.n1337 147.374
R2196 VSS.n1335 VSS.n1334 147.374
R2197 VSS.n1330 VSS.n1284 147.374
R2198 VSS.n1328 VSS.n1327 147.374
R2199 VSS.n1323 VSS.n1287 147.374
R2200 VSS.n1321 VSS.n1320 147.374
R2201 VSS.n1316 VSS.n1290 147.374
R2202 VSS.n1314 VSS.n1313 147.374
R2203 VSS.n1309 VSS.n1293 147.374
R2204 VSS.n1307 VSS.n1306 147.374
R2205 VSS.n1302 VSS.n1301 147.374
R2206 VSS.n1638 VSS.n509 147.374
R2207 VSS.n524 VSS.n514 147.374
R2208 VSS.n528 VSS.n515 147.374
R2209 VSS.n532 VSS.n516 147.374
R2210 VSS.n536 VSS.n517 147.374
R2211 VSS.n540 VSS.n518 147.374
R2212 VSS.n544 VSS.n519 147.374
R2213 VSS.n548 VSS.n520 147.374
R2214 VSS.n552 VSS.n521 147.374
R2215 VSS.n556 VSS.n522 147.374
R2216 VSS.n562 VSS.n561 147.374
R2217 VSS.n2140 VSS.n2139 147.374
R2218 VSS.n2137 VSS.n2132 147.374
R2219 VSS.n2314 VSS.n2313 147.374
R2220 VSS.n145 VSS.n143 147.374
R2221 VSS.n2138 VSS.n2137 147.374
R2222 VSS.n2141 VSS.n2140 147.374
R2223 VSS.n2313 VSS.n141 147.374
R2224 VSS.n2307 VSS.n143 147.374
R2225 VSS.n1639 VSS.n1638 147.374
R2226 VSS.n527 VSS.n514 147.374
R2227 VSS.n531 VSS.n515 147.374
R2228 VSS.n535 VSS.n516 147.374
R2229 VSS.n539 VSS.n517 147.374
R2230 VSS.n543 VSS.n518 147.374
R2231 VSS.n547 VSS.n519 147.374
R2232 VSS.n551 VSS.n520 147.374
R2233 VSS.n555 VSS.n521 147.374
R2234 VSS.n523 VSS.n522 147.374
R2235 VSS.n562 VSS.n506 147.374
R2236 VSS.n1301 VSS.n1294 147.374
R2237 VSS.n1308 VSS.n1307 147.374
R2238 VSS.n1293 VSS.n1291 147.374
R2239 VSS.n1315 VSS.n1314 147.374
R2240 VSS.n1290 VSS.n1288 147.374
R2241 VSS.n1322 VSS.n1321 147.374
R2242 VSS.n1287 VSS.n1285 147.374
R2243 VSS.n1329 VSS.n1328 147.374
R2244 VSS.n1284 VSS.n1282 147.374
R2245 VSS.n1336 VSS.n1335 147.374
R2246 VSS.n1339 VSS.n1338 147.374
R2247 VSS.n1594 VSS.n607 147.374
R2248 VSS.n1588 VSS.n609 147.374
R2249 VSS.n1584 VSS.n610 147.374
R2250 VSS.n1580 VSS.n611 147.374
R2251 VSS.n1576 VSS.n612 147.374
R2252 VSS.n1572 VSS.n613 147.374
R2253 VSS.n1568 VSS.n614 147.374
R2254 VSS.n1564 VSS.n615 147.374
R2255 VSS.n1560 VSS.n616 147.374
R2256 VSS.n1556 VSS.n617 147.374
R2257 VSS.n1552 VSS.n618 147.374
R2258 VSS.n986 VSS.n985 147.374
R2259 VSS.n981 VSS.n935 147.374
R2260 VSS.n979 VSS.n978 147.374
R2261 VSS.n974 VSS.n973 147.374
R2262 VSS.n971 VSS.n970 147.374
R2263 VSS.n966 VSS.n965 147.374
R2264 VSS.n963 VSS.n962 147.374
R2265 VSS.n958 VSS.n957 147.374
R2266 VSS.n955 VSS.n954 147.374
R2267 VSS.n950 VSS.n949 147.374
R2268 VSS.n947 VSS.n946 147.374
R2269 VSS.n2623 VSS.n36 147.374
R2270 VSS.n2615 VSS.n22 147.374
R2271 VSS.n2611 VSS.n23 147.374
R2272 VSS.n2606 VSS.n24 147.374
R2273 VSS.n27 VSS.n25 147.374
R2274 VSS.n30 VSS.n19 147.374
R2275 VSS.n2625 VSS.n20 147.374
R2276 VSS.n2583 VSS.n31 147.374
R2277 VSS.n2587 VSS.n32 147.374
R2278 VSS.n2591 VSS.n33 147.374
R2279 VSS.n2594 VSS.n34 147.374
R2280 VSS.n1499 VSS.n625 147.374
R2281 VSS.n1503 VSS.n626 147.374
R2282 VSS.n1507 VSS.n627 147.374
R2283 VSS.n1511 VSS.n628 147.374
R2284 VSS.n1515 VSS.n629 147.374
R2285 VSS.n1519 VSS.n630 147.374
R2286 VSS.n1523 VSS.n631 147.374
R2287 VSS.n1527 VSS.n632 147.374
R2288 VSS.n1531 VSS.n633 147.374
R2289 VSS.n1535 VSS.n634 147.374
R2290 VSS.n637 VSS.n635 147.374
R2291 VSS.n1999 VSS.n1998 147.374
R2292 VSS.n1993 VSS.n344 147.374
R2293 VSS.n1991 VSS.n1990 147.374
R2294 VSS.n1986 VSS.n1985 147.374
R2295 VSS.n1983 VSS.n1982 147.374
R2296 VSS.n1978 VSS.n1977 147.374
R2297 VSS.n1975 VSS.n1974 147.374
R2298 VSS.n1968 VSS.n1967 147.374
R2299 VSS.n1963 VSS.n354 147.374
R2300 VSS.n1952 VSS.n356 147.374
R2301 VSS.n1955 VSS.n1954 147.374
R2302 VSS.n1948 VSS.n362 147.374
R2303 VSS.n1946 VSS.n1945 147.374
R2304 VSS.n1941 VSS.n1940 147.374
R2305 VSS.n1938 VSS.n1937 147.374
R2306 VSS.n1933 VSS.n1932 147.374
R2307 VSS.n1930 VSS.n1929 147.374
R2308 VSS.n1925 VSS.n1924 147.374
R2309 VSS.n1922 VSS.n1921 147.374
R2310 VSS.n1831 VSS.n379 147.374
R2311 VSS.n1757 VSS.n380 147.374
R2312 VSS.n1761 VSS.n381 147.374
R2313 VSS.n1765 VSS.n382 147.374
R2314 VSS.n1769 VSS.n383 147.374
R2315 VSS.n1773 VSS.n384 147.374
R2316 VSS.n1777 VSS.n385 147.374
R2317 VSS.n1781 VSS.n386 147.374
R2318 VSS.n406 VSS.n387 147.374
R2319 VSS.n1789 VSS.n388 147.374
R2320 VSS.n1793 VSS.n389 147.374
R2321 VSS.n1800 VSS.n390 147.374
R2322 VSS.n1804 VSS.n391 147.374
R2323 VSS.n1808 VSS.n392 147.374
R2324 VSS.n1812 VSS.n393 147.374
R2325 VSS.n1816 VSS.n394 147.374
R2326 VSS.n1820 VSS.n395 147.374
R2327 VSS.n1824 VSS.n396 147.374
R2328 VSS.n398 VSS.n397 147.374
R2329 VSS.n2397 VSS.n2396 147.374
R2330 VSS.n2391 VSS.n106 147.374
R2331 VSS.n2388 VSS.n107 147.374
R2332 VSS.n2384 VSS.n108 147.374
R2333 VSS.n2380 VSS.n109 147.374
R2334 VSS.n2376 VSS.n110 147.374
R2335 VSS.n2372 VSS.n111 147.374
R2336 VSS.n2368 VSS.n112 147.374
R2337 VSS.n2364 VSS.n113 147.374
R2338 VSS.n2401 VSS.n2400 147.374
R2339 VSS.n2407 VSS.n2406 147.374
R2340 VSS.n2410 VSS.n2409 147.374
R2341 VSS.n2415 VSS.n2414 147.374
R2342 VSS.n2418 VSS.n2417 147.374
R2343 VSS.n2423 VSS.n2422 147.374
R2344 VSS.n2426 VSS.n2425 147.374
R2345 VSS.n2431 VSS.n2430 147.374
R2346 VSS.n2434 VSS.n2433 147.374
R2347 VSS.n2439 VSS.n2438 147.374
R2348 VSS.n2442 VSS.n2441 147.374
R2349 VSS.n2447 VSS.n2446 147.374
R2350 VSS.n2450 VSS.n2449 147.374
R2351 VSS.n2455 VSS.n2454 147.374
R2352 VSS.n2458 VSS.n2457 147.374
R2353 VSS.n2463 VSS.n2462 147.374
R2354 VSS.n2466 VSS.n2465 147.374
R2355 VSS.n2471 VSS.n2470 147.374
R2356 VSS.n2474 VSS.n2473 147.374
R2357 VSS.n2479 VSS.n2478 147.374
R2358 VSS.n2482 VSS.n2481 147.374
R2359 VSS.n2487 VSS.n2486 147.374
R2360 VSS.n2490 VSS.n2489 147.374
R2361 VSS.n2495 VSS.n2494 147.374
R2362 VSS.n2498 VSS.n2497 147.374
R2363 VSS.n2503 VSS.n2502 147.374
R2364 VSS.n2506 VSS.n2505 147.374
R2365 VSS.n2511 VSS.n2510 147.374
R2366 VSS.n2514 VSS.n2513 147.374
R2367 VSS.n2519 VSS.n2518 147.374
R2368 VSS.n2522 VSS.n2521 147.374
R2369 VSS.n2527 VSS.n2526 147.374
R2370 VSS.n2530 VSS.n2529 147.374
R2371 VSS.n2535 VSS.n2534 147.374
R2372 VSS.n2538 VSS.n2537 147.374
R2373 VSS.n2543 VSS.n2542 147.374
R2374 VSS.n1092 VSS.n769 147.374
R2375 VSS.n1099 VSS.n1098 147.374
R2376 VSS.n1100 VSS.n767 147.374
R2377 VSS.n1107 VSS.n1106 147.374
R2378 VSS.n1108 VSS.n765 147.374
R2379 VSS.n1115 VSS.n1114 147.374
R2380 VSS.n1116 VSS.n763 147.374
R2381 VSS.n1123 VSS.n1122 147.374
R2382 VSS.n1124 VSS.n761 147.374
R2383 VSS.n1131 VSS.n1130 147.374
R2384 VSS.n1132 VSS.n724 147.374
R2385 VSS.n1140 VSS.n726 147.374
R2386 VSS.n1144 VSS.n727 147.374
R2387 VSS.n1148 VSS.n728 147.374
R2388 VSS.n1152 VSS.n729 147.374
R2389 VSS.n1156 VSS.n730 147.374
R2390 VSS.n1160 VSS.n731 147.374
R2391 VSS.n1164 VSS.n732 147.374
R2392 VSS.n1168 VSS.n733 147.374
R2393 VSS.n1172 VSS.n734 147.374
R2394 VSS.n1176 VSS.n735 147.374
R2395 VSS.n1180 VSS.n736 147.374
R2396 VSS.n1188 VSS.n738 147.374
R2397 VSS.n1192 VSS.n739 147.374
R2398 VSS.n1196 VSS.n740 147.374
R2399 VSS.n1200 VSS.n741 147.374
R2400 VSS.n1204 VSS.n742 147.374
R2401 VSS.n1208 VSS.n743 147.374
R2402 VSS.n1212 VSS.n744 147.374
R2403 VSS.n1216 VSS.n745 147.374
R2404 VSS.n1220 VSS.n746 147.374
R2405 VSS.n1224 VSS.n747 147.374
R2406 VSS.n1228 VSS.n748 147.374
R2407 VSS.n1236 VSS.n750 147.374
R2408 VSS.n1240 VSS.n751 147.374
R2409 VSS.n1244 VSS.n752 147.374
R2410 VSS.n1248 VSS.n753 147.374
R2411 VSS.n1252 VSS.n754 147.374
R2412 VSS.n1256 VSS.n755 147.374
R2413 VSS.n1260 VSS.n756 147.374
R2414 VSS.n1264 VSS.n757 147.374
R2415 VSS.n1268 VSS.n758 147.374
R2416 VSS.n1275 VSS.n759 147.374
R2417 VSS.n1346 VSS.n722 147.374
R2418 VSS.n1347 VSS.n1346 147.374
R2419 VSS.n1275 VSS.n1274 147.374
R2420 VSS.n1270 VSS.n758 147.374
R2421 VSS.n1267 VSS.n757 147.374
R2422 VSS.n1263 VSS.n756 147.374
R2423 VSS.n1259 VSS.n755 147.374
R2424 VSS.n1255 VSS.n754 147.374
R2425 VSS.n1251 VSS.n753 147.374
R2426 VSS.n1247 VSS.n752 147.374
R2427 VSS.n1243 VSS.n751 147.374
R2428 VSS.n1239 VSS.n750 147.374
R2429 VSS.n1231 VSS.n748 147.374
R2430 VSS.n1227 VSS.n747 147.374
R2431 VSS.n1223 VSS.n746 147.374
R2432 VSS.n1219 VSS.n745 147.374
R2433 VSS.n1215 VSS.n744 147.374
R2434 VSS.n1211 VSS.n743 147.374
R2435 VSS.n1207 VSS.n742 147.374
R2436 VSS.n1203 VSS.n741 147.374
R2437 VSS.n1199 VSS.n740 147.374
R2438 VSS.n1195 VSS.n739 147.374
R2439 VSS.n1191 VSS.n738 147.374
R2440 VSS.n1183 VSS.n736 147.374
R2441 VSS.n1179 VSS.n735 147.374
R2442 VSS.n1175 VSS.n734 147.374
R2443 VSS.n1171 VSS.n733 147.374
R2444 VSS.n1167 VSS.n732 147.374
R2445 VSS.n1163 VSS.n731 147.374
R2446 VSS.n1159 VSS.n730 147.374
R2447 VSS.n1155 VSS.n729 147.374
R2448 VSS.n1151 VSS.n728 147.374
R2449 VSS.n1147 VSS.n727 147.374
R2450 VSS.n1143 VSS.n726 147.374
R2451 VSS.n1135 VSS.n724 147.374
R2452 VSS.n1130 VSS.n1129 147.374
R2453 VSS.n1125 VSS.n1124 147.374
R2454 VSS.n1122 VSS.n1121 147.374
R2455 VSS.n1117 VSS.n1116 147.374
R2456 VSS.n1114 VSS.n1113 147.374
R2457 VSS.n1109 VSS.n1108 147.374
R2458 VSS.n1106 VSS.n1105 147.374
R2459 VSS.n1101 VSS.n1100 147.374
R2460 VSS.n1098 VSS.n1097 147.374
R2461 VSS.n1093 VSS.n1092 147.374
R2462 VSS.n2397 VSS.n115 147.374
R2463 VSS.n2389 VSS.n106 147.374
R2464 VSS.n2385 VSS.n107 147.374
R2465 VSS.n2381 VSS.n108 147.374
R2466 VSS.n2377 VSS.n109 147.374
R2467 VSS.n2373 VSS.n110 147.374
R2468 VSS.n2369 VSS.n111 147.374
R2469 VSS.n2365 VSS.n112 147.374
R2470 VSS.n113 VSS.n103 147.374
R2471 VSS.n2402 VSS.n2401 147.374
R2472 VSS.n2408 VSS.n2407 147.374
R2473 VSS.n2409 VSS.n99 147.374
R2474 VSS.n2416 VSS.n2415 147.374
R2475 VSS.n2417 VSS.n97 147.374
R2476 VSS.n2424 VSS.n2423 147.374
R2477 VSS.n2425 VSS.n95 147.374
R2478 VSS.n2432 VSS.n2431 147.374
R2479 VSS.n2433 VSS.n93 147.374
R2480 VSS.n2440 VSS.n2439 147.374
R2481 VSS.n2441 VSS.n91 147.374
R2482 VSS.n2448 VSS.n2447 147.374
R2483 VSS.n2449 VSS.n89 147.374
R2484 VSS.n2456 VSS.n2455 147.374
R2485 VSS.n2457 VSS.n87 147.374
R2486 VSS.n2464 VSS.n2463 147.374
R2487 VSS.n2465 VSS.n85 147.374
R2488 VSS.n2472 VSS.n2471 147.374
R2489 VSS.n2473 VSS.n83 147.374
R2490 VSS.n2480 VSS.n2479 147.374
R2491 VSS.n2481 VSS.n81 147.374
R2492 VSS.n2488 VSS.n2487 147.374
R2493 VSS.n2489 VSS.n79 147.374
R2494 VSS.n2496 VSS.n2495 147.374
R2495 VSS.n2497 VSS.n77 147.374
R2496 VSS.n2504 VSS.n2503 147.374
R2497 VSS.n2505 VSS.n75 147.374
R2498 VSS.n2512 VSS.n2511 147.374
R2499 VSS.n2513 VSS.n73 147.374
R2500 VSS.n2520 VSS.n2519 147.374
R2501 VSS.n2521 VSS.n71 147.374
R2502 VSS.n2528 VSS.n2527 147.374
R2503 VSS.n2529 VSS.n69 147.374
R2504 VSS.n2536 VSS.n2535 147.374
R2505 VSS.n2537 VSS.n67 147.374
R2506 VSS.n2544 VSS.n2543 147.374
R2507 VSS.n672 VSS.n666 140.69
R2508 VSS.n673 VSS.n672 140.69
R2509 VSS.n673 VSS.n662 140.69
R2510 VSS.n680 VSS.n662 140.69
R2511 VSS.n681 VSS.n680 140.69
R2512 VSS.n681 VSS.n658 140.69
R2513 VSS.n688 VSS.n658 140.69
R2514 VSS.n1466 VSS.n1434 140.69
R2515 VSS.n1459 VSS.n1434 140.69
R2516 VSS.n1459 VSS.n1458 140.69
R2517 VSS.n1458 VSS.n1438 140.69
R2518 VSS.n1451 VSS.n1438 140.69
R2519 VSS.n1451 VSS.n1450 140.69
R2520 VSS.n1450 VSS.n1442 140.69
R2521 VSS.n825 VSS.n824 140.69
R2522 VSS.n824 VSS.n798 140.69
R2523 VSS.n817 VSS.n798 140.69
R2524 VSS.n817 VSS.n816 140.69
R2525 VSS.n816 VSS.n802 140.69
R2526 VSS.n809 VSS.n802 140.69
R2527 VSS.n809 VSS.n808 140.69
R2528 VSS.n852 VSS.n847 140.69
R2529 VSS.n859 VSS.n847 140.69
R2530 VSS.n860 VSS.n859 140.69
R2531 VSS.n860 VSS.n843 140.69
R2532 VSS.n868 VSS.n843 140.69
R2533 VSS.n869 VSS.n868 140.69
R2534 VSS.n869 VSS.n840 140.69
R2535 VSS.n476 VSS.n452 140.69
R2536 VSS.n469 VSS.n452 140.69
R2537 VSS.n423 VSS.n422 140.69
R2538 VSS.n423 VSS.n414 140.69
R2539 VSS.n2231 VSS.n198 117.233
R2540 VSS.n2146 VSS.n2129 99.5348
R2541 VSS.n2152 VSS.n2129 99.5348
R2542 VSS.n2152 VSS.n2125 99.5348
R2543 VSS.n2158 VSS.n2125 99.5348
R2544 VSS.n2158 VSS.n2121 99.5348
R2545 VSS.n2165 VSS.n2121 99.5348
R2546 VSS.n2165 VSS.n2164 99.5348
R2547 VSS.n2171 VSS.n235 99.5348
R2548 VSS.n2177 VSS.n235 99.5348
R2549 VSS.n2177 VSS.n231 99.5348
R2550 VSS.n2183 VSS.n231 99.5348
R2551 VSS.n2183 VSS.n227 99.5348
R2552 VSS.n2189 VSS.n227 99.5348
R2553 VSS.n2189 VSS.n223 99.5348
R2554 VSS.n2195 VSS.n223 99.5348
R2555 VSS.n2195 VSS.n219 99.5348
R2556 VSS.n2201 VSS.n219 99.5348
R2557 VSS.n2201 VSS.n215 99.5348
R2558 VSS.n2207 VSS.n215 99.5348
R2559 VSS.n2207 VSS.n211 99.5348
R2560 VSS.n2213 VSS.n211 99.5348
R2561 VSS.n2213 VSS.n207 99.5348
R2562 VSS.n2219 VSS.n207 99.5348
R2563 VSS.n2219 VSS.n203 99.5348
R2564 VSS.n2225 VSS.n203 99.5348
R2565 VSS.n1090 VSS.n1089 99.5348
R2566 VSS.n1088 VSS.n772 99.5348
R2567 VSS.n901 VSS.n772 99.5348
R2568 VSS.n904 VSS.n901 99.5348
R2569 VSS.n912 VSS.n896 99.5348
R2570 VSS.n913 VSS.n912 99.5348
R2571 VSS.n914 VSS.n913 99.5348
R2572 VSS.n916 VSS.n892 99.5348
R2573 VSS.n922 VSS.n892 99.5348
R2574 VSS.n923 VSS.n922 99.5348
R2575 VSS.n924 VSS.n887 99.5348
R2576 VSS.n933 VSS.n887 99.5348
R2577 VSS.n1073 VSS.n1071 99.5348
R2578 VSS.n1073 VSS.n1072 99.5348
R2579 VSS.n1022 VSS.n1020 99.5348
R2580 VSS.n1022 VSS.n1021 99.5348
R2581 VSS.n1021 VSS.n1002 99.5348
R2582 VSS.n1048 VSS.n1003 99.5348
R2583 VSS.n1042 VSS.n1003 99.5348
R2584 VSS.n1042 VSS.n1041 99.5348
R2585 VSS.n1038 VSS.n1037 99.5348
R2586 VSS.n1037 VSS.n1036 99.5348
R2587 VSS.n1036 VSS.n1010 99.5348
R2588 VSS.n2353 VSS.n123 99.5348
R2589 VSS.n2354 VSS.n2353 99.5348
R2590 VSS.n2355 VSS.n2354 99.5348
R2591 VSS.n121 VSS.n105 99.5348
R2592 VSS.n1089 VSS.t30 92.2161
R2593 VSS.n121 VSS.t2 92.2161
R2594 VSS.n1680 VSS.t86 90.6265
R2595 VSS.n1664 VSS.t79 90.6265
R2596 VSS.n1736 VSS.t96 90.6265
R2597 VSS.n1719 VSS.t89 90.6265
R2598 VSS.n1071 VSS.t33 89.2886
R2599 VSS.n1072 VSS.t22 89.2886
R2600 VSS.n2144 VSS.n2143 85.8358
R2601 VSS.n2148 VSS.n2131 85.8358
R2602 VSS.n2308 VSS.n147 85.8358
R2603 VSS.n1539 VSS.n638 82.4476
R2604 VSS.n2621 VSS.n2602 82.4476
R2605 VSS.n1497 VSS.n639 82.4476
R2606 VSS.n2596 VSS.n2595 82.4476
R2607 VSS.n1626 VSS.n574 82.4476
R2608 VSS.n989 VSS.n988 82.4476
R2609 VSS.n1597 VSS.n1596 82.4476
R2610 VSS.n1553 VSS.n620 82.4476
R2611 VSS.n1342 VSS.n1341 82.4476
R2612 VSS.n1642 VSS.n1641 82.4476
R2613 VSS.n1303 VSS.n1300 82.4476
R2614 VSS.n454 VSS.t90 81.8918
R2615 VSS.n467 VSS.t114 81.8918
R2616 VSS.n413 VSS.t125 81.8918
R2617 VSS.n430 VSS.t123 81.8918
R2618 VSS.n1680 VSS.t84 81.8918
R2619 VSS.n1679 VSS.t127 81.8918
R2620 VSS.n1664 VSS.t76 81.8918
R2621 VSS.n1740 VSS.t93 81.8918
R2622 VSS.n1736 VSS.t95 81.8918
R2623 VSS.n1719 VSS.t87 81.8918
R2624 VSS.n1069 VSS.n933 79.0424
R2625 VSS.n1828 VSS.n374 76.8005
R2626 VSS.n2002 VSS.n2001 76.8005
R2627 VSS.n1920 VSS.n1919 76.8005
R2628 VSS.n1834 VSS.n1833 76.8005
R2629 VSS.n1094 VSS.n770 76.8005
R2630 VSS.n1349 VSS.n1348 76.8005
R2631 VSS.n2395 VSS.n2361 76.8005
R2632 VSS.n2549 VSS.n64 76.8005
R2633 VSS.n2164 VSS.n2117 74.6512
R2634 VSS.n904 VSS.t43 71.7237
R2635 VSS.t60 VSS.n123 71.7237
R2636 VSS.t73 VSS.n666 70.3453
R2637 VSS.t75 VSS.n1466 70.3453
R2638 VSS.n808 VSS.t111 70.3453
R2639 VSS.t68 VSS.n840 70.3453
R2640 VSS.n469 VSS.t116 70.3453
R2641 VSS.t126 VSS.n414 70.3453
R2642 VSS.n924 VSS.t8 68.7962
R2643 VSS.t11 VSS.n1002 68.7962
R2644 VSS.n2624 VSS.n21 66.162
R2645 VSS.n1138 VSS.n1137 64.7534
R2646 VSS.n2405 VSS.n2404 64.7534
R2647 VSS.n2316 VSS.n138 62.1181
R2648 VSS.n1345 VSS.n723 61.9943
R2649 VSS.n1830 VSS.n376 54.18
R2650 VSS.n2004 VSS.n341 54.18
R2651 VSS.n914 VSS.t9 51.2314
R2652 VSS.n1038 VSS.t10 51.2314
R2653 VSS.n2225 VSS.t49 49.7676
R2654 VSS.n916 VSS.t9 48.3039
R2655 VSS.n1041 VSS.t10 48.3039
R2656 VSS.n559 VSS.n503 45.3391
R2657 VSS.n1186 VSS.n1185 39.1534
R2658 VSS.n1234 VSS.n1233 39.1534
R2659 VSS.n2453 VSS.n2452 39.1534
R2660 VSS.n2501 VSS.n2500 39.1534
R2661 VSS.t49 VSS.n198 38.2032
R2662 VSS.n1839 VSS.n376 35.4256
R2663 VSS.n1839 VSS.n1838 35.4256
R2664 VSS.n1845 VSS.n239 35.4256
R2665 VSS.n2110 VSS.n246 35.4256
R2666 VSS.n2110 VSS.n2109 35.4256
R2667 VSS.n2109 VSS.n2108 35.4256
R2668 VSS.n2102 VSS.n253 35.4256
R2669 VSS.n2102 VSS.n2101 35.4256
R2670 VSS.n2101 VSS.n2100 35.4256
R2671 VSS.n2094 VSS.n260 35.4256
R2672 VSS.n2094 VSS.n2093 35.4256
R2673 VSS.n2093 VSS.n2092 35.4256
R2674 VSS.n2086 VSS.n267 35.4256
R2675 VSS.n2086 VSS.n2085 35.4256
R2676 VSS.n2085 VSS.n2084 35.4256
R2677 VSS.n2078 VSS.n274 35.4256
R2678 VSS.n2078 VSS.n2077 35.4256
R2679 VSS.n2076 VSS.n278 35.4256
R2680 VSS.n2070 VSS.n278 35.4256
R2681 VSS.n2070 VSS.n2069 35.4256
R2682 VSS.n2068 VSS.n285 35.4256
R2683 VSS.n2062 VSS.n285 35.4256
R2684 VSS.n2062 VSS.n2061 35.4256
R2685 VSS.n2060 VSS.n292 35.4256
R2686 VSS.n2054 VSS.n292 35.4256
R2687 VSS.n2054 VSS.n2053 35.4256
R2688 VSS.n2052 VSS.n299 35.4256
R2689 VSS.n2046 VSS.n299 35.4256
R2690 VSS.n2045 VSS.n2044 35.4256
R2691 VSS.n2044 VSS.n306 35.4256
R2692 VSS.n2038 VSS.n306 35.4256
R2693 VSS.n2037 VSS.n2036 35.4256
R2694 VSS.n2036 VSS.n313 35.4256
R2695 VSS.n2030 VSS.n313 35.4256
R2696 VSS.n2029 VSS.n2028 35.4256
R2697 VSS.n2028 VSS.n320 35.4256
R2698 VSS.n2022 VSS.n320 35.4256
R2699 VSS.n2021 VSS.n2020 35.4256
R2700 VSS.n2020 VSS.n327 35.4256
R2701 VSS.n2014 VSS.n327 35.4256
R2702 VSS.n2013 VSS.n2012 35.4256
R2703 VSS.n2012 VSS.n334 35.4256
R2704 VSS.n2006 VSS.n2005 35.4256
R2705 VSS.n2005 VSS.n2004 35.4256
R2706 VSS.n1344 VSS.n1278 35.4256
R2707 VSS.n1383 VSS.n513 35.4256
R2708 VSS.n1636 VSS.n563 35.4256
R2709 VSS.n1630 VSS.n1629 35.4256
R2710 VSS.n1549 VSS.n608 35.4256
R2711 VSS.n1543 VSS.n1542 35.4256
R2712 VSS.n645 VSS.n624 35.4256
R2713 VSS.n2569 VSS.n44 35.4256
R2714 VSS.n2575 VSS.n44 35.4256
R2715 VSS.n2575 VSS.n45 35.4256
R2716 VSS.n2599 VSS.n21 35.4256
R2717 VSS.n274 VSS.t53 34.9046
R2718 VSS.n2046 VSS.t24 34.9046
R2719 VSS.n1845 VSS.t88 33.8627
R2720 VSS.t77 VSS.n334 33.8627
R2721 VSS.n1671 VSS.n1670 32.8962
R2722 VSS.n1726 VSS.n1725 32.8962
R2723 VSS.t8 VSS.n923 30.739
R2724 VSS.t11 VSS.n1048 30.739
R2725 VSS.n2117 VSS.n2116 30.7369
R2726 VSS.n2116 VSS.t36 29.695
R2727 VSS.t91 VSS.n2013 29.695
R2728 VSS.n2077 VSS.t55 28.6531
R2729 VSS.t3 VSS.n2052 28.6531
R2730 VSS.n470 VSS.n468 28.3989
R2731 VSS.n427 VSS.n426 28.3989
R2732 VSS.n1695 VSS.n1694 27.9576
R2733 VSS.n1699 VSS.n1698 27.9576
R2734 VSS.n1703 VSS.n1702 27.9576
R2735 VSS.n1707 VSS.n1706 27.9576
R2736 VSS.n1711 VSS.n1710 27.9576
R2737 VSS.t43 VSS.n896 27.8115
R2738 VSS.n1010 VSS.t60 27.8115
R2739 VSS.n1693 VSS.n1692 27.7293
R2740 VSS.n1697 VSS.n1696 27.7293
R2741 VSS.n1701 VSS.n1700 27.7293
R2742 VSS.n1705 VSS.n1704 27.7293
R2743 VSS.n1709 VSS.n1708 27.7293
R2744 VSS.n1713 VSS.n1712 27.7293
R2745 VSS.n448 VSS.n447 27.7293
R2746 VSS.n446 VSS.n445 27.7293
R2747 VSS.n444 VSS.n443 27.7293
R2748 VSS.n442 VSS.n441 27.7293
R2749 VSS.n440 VSS.n439 27.7293
R2750 VSS.n267 VSS.t16 27.6112
R2751 VSS.n2038 VSS.t20 27.6112
R2752 VSS.n1542 VSS.n1541 27.6112
R2753 VSS.n464 VSS.n455 27.5286
R2754 VSS.n435 VSS.n412 27.5286
R2755 VSS.n1687 VSS.n1658 27.5286
R2756 VSS.n1688 VSS.n1656 27.5286
R2757 VSS.n1748 VSS.n1731 27.5286
R2758 VSS.n1747 VSS.n1733 27.5286
R2759 VSS.n690 VSS.n689 25.6009
R2760 VSS.n1444 VSS.n694 25.6009
R2761 VSS.n829 VSS.n795 25.6009
R2762 VSS.n851 VSS.n839 25.6009
R2763 VSS.n638 VSS.n54 25.6005
R2764 VSS.n2559 VSS.n54 25.6005
R2765 VSS.n2560 VSS.n2559 25.6005
R2766 VSS.n2561 VSS.n2560 25.6005
R2767 VSS.n2561 VSS.n47 25.6005
R2768 VSS.n2571 VSS.n47 25.6005
R2769 VSS.n2572 VSS.n2571 25.6005
R2770 VSS.n2573 VSS.n2572 25.6005
R2771 VSS.n2573 VSS.n38 25.6005
R2772 VSS.n2601 VSS.n38 25.6005
R2773 VSS.n2602 VSS.n2601 25.6005
R2774 VSS.n1539 VSS.n1538 25.6005
R2775 VSS.n1538 VSS.n1537 25.6005
R2776 VSS.n1537 VSS.n1534 25.6005
R2777 VSS.n1534 VSS.n1533 25.6005
R2778 VSS.n1533 VSS.n1530 25.6005
R2779 VSS.n1530 VSS.n1529 25.6005
R2780 VSS.n1529 VSS.n1526 25.6005
R2781 VSS.n1526 VSS.n1525 25.6005
R2782 VSS.n1525 VSS.n1522 25.6005
R2783 VSS.n1522 VSS.n1521 25.6005
R2784 VSS.n1521 VSS.n1518 25.6005
R2785 VSS.n1518 VSS.n1517 25.6005
R2786 VSS.n1517 VSS.n1514 25.6005
R2787 VSS.n1514 VSS.n1513 25.6005
R2788 VSS.n1513 VSS.n1510 25.6005
R2789 VSS.n1510 VSS.n1509 25.6005
R2790 VSS.n1509 VSS.n1506 25.6005
R2791 VSS.n1506 VSS.n1505 25.6005
R2792 VSS.n1505 VSS.n1502 25.6005
R2793 VSS.n1502 VSS.n1501 25.6005
R2794 VSS.n1501 VSS.n1498 25.6005
R2795 VSS.n1498 VSS.n1497 25.6005
R2796 VSS.n641 VSS.n639 25.6005
R2797 VSS.n641 VSS.n640 25.6005
R2798 VSS.n640 VSS.n50 25.6005
R2799 VSS.n2565 VSS.n50 25.6005
R2800 VSS.n2566 VSS.n2565 25.6005
R2801 VSS.n2567 VSS.n2566 25.6005
R2802 VSS.n2567 VSS.n42 25.6005
R2803 VSS.n2577 VSS.n42 25.6005
R2804 VSS.n2578 VSS.n2577 25.6005
R2805 VSS.n2597 VSS.n2578 25.6005
R2806 VSS.n2597 VSS.n2596 25.6005
R2807 VSS.n2621 VSS.n2620 25.6005
R2808 VSS.n2620 VSS.n2619 25.6005
R2809 VSS.n2619 VSS.n2618 25.6005
R2810 VSS.n2618 VSS.n2616 25.6005
R2811 VSS.n2616 VSS.n2613 25.6005
R2812 VSS.n2613 VSS.n2612 25.6005
R2813 VSS.n2607 VSS.n2604 25.6005
R2814 VSS.n28 VSS.n18 25.6005
R2815 VSS.n2581 VSS.n2579 25.6005
R2816 VSS.n2582 VSS.n2581 25.6005
R2817 VSS.n2585 VSS.n2582 25.6005
R2818 VSS.n2586 VSS.n2585 25.6005
R2819 VSS.n2589 VSS.n2586 25.6005
R2820 VSS.n2590 VSS.n2589 25.6005
R2821 VSS.n2593 VSS.n2590 25.6005
R2822 VSS.n2595 VSS.n2593 25.6005
R2823 VSS.n1841 VSS.n374 25.6005
R2824 VSS.n1842 VSS.n1841 25.6005
R2825 VSS.n1843 VSS.n1842 25.6005
R2826 VSS.n1843 VSS.n243 25.6005
R2827 VSS.n2114 VSS.n243 25.6005
R2828 VSS.n2114 VSS.n2113 25.6005
R2829 VSS.n2113 VSS.n2112 25.6005
R2830 VSS.n2112 VSS.n244 25.6005
R2831 VSS.n2106 VSS.n244 25.6005
R2832 VSS.n2106 VSS.n2105 25.6005
R2833 VSS.n2105 VSS.n2104 25.6005
R2834 VSS.n2104 VSS.n251 25.6005
R2835 VSS.n2098 VSS.n251 25.6005
R2836 VSS.n2098 VSS.n2097 25.6005
R2837 VSS.n2097 VSS.n2096 25.6005
R2838 VSS.n2096 VSS.n258 25.6005
R2839 VSS.n2090 VSS.n258 25.6005
R2840 VSS.n2090 VSS.n2089 25.6005
R2841 VSS.n2089 VSS.n2088 25.6005
R2842 VSS.n2088 VSS.n265 25.6005
R2843 VSS.n2082 VSS.n265 25.6005
R2844 VSS.n2082 VSS.n2081 25.6005
R2845 VSS.n2081 VSS.n2080 25.6005
R2846 VSS.n2080 VSS.n272 25.6005
R2847 VSS.n2074 VSS.n272 25.6005
R2848 VSS.n2074 VSS.n2073 25.6005
R2849 VSS.n2073 VSS.n2072 25.6005
R2850 VSS.n2072 VSS.n280 25.6005
R2851 VSS.n2066 VSS.n280 25.6005
R2852 VSS.n2066 VSS.n2065 25.6005
R2853 VSS.n2065 VSS.n2064 25.6005
R2854 VSS.n2064 VSS.n287 25.6005
R2855 VSS.n2058 VSS.n287 25.6005
R2856 VSS.n2058 VSS.n2057 25.6005
R2857 VSS.n2057 VSS.n2056 25.6005
R2858 VSS.n2056 VSS.n294 25.6005
R2859 VSS.n2050 VSS.n294 25.6005
R2860 VSS.n2050 VSS.n2049 25.6005
R2861 VSS.n2049 VSS.n2048 25.6005
R2862 VSS.n2048 VSS.n301 25.6005
R2863 VSS.n2042 VSS.n301 25.6005
R2864 VSS.n2042 VSS.n2041 25.6005
R2865 VSS.n2041 VSS.n2040 25.6005
R2866 VSS.n2040 VSS.n308 25.6005
R2867 VSS.n2034 VSS.n308 25.6005
R2868 VSS.n2034 VSS.n2033 25.6005
R2869 VSS.n2033 VSS.n2032 25.6005
R2870 VSS.n2032 VSS.n315 25.6005
R2871 VSS.n2026 VSS.n315 25.6005
R2872 VSS.n2026 VSS.n2025 25.6005
R2873 VSS.n2025 VSS.n2024 25.6005
R2874 VSS.n2024 VSS.n322 25.6005
R2875 VSS.n2018 VSS.n322 25.6005
R2876 VSS.n2018 VSS.n2017 25.6005
R2877 VSS.n2017 VSS.n2016 25.6005
R2878 VSS.n2016 VSS.n329 25.6005
R2879 VSS.n2010 VSS.n329 25.6005
R2880 VSS.n2010 VSS.n2009 25.6005
R2881 VSS.n2009 VSS.n2008 25.6005
R2882 VSS.n2008 VSS.n336 25.6005
R2883 VSS.n2002 VSS.n336 25.6005
R2884 VSS.n2001 VSS.n2000 25.6005
R2885 VSS.n2000 VSS.n343 25.6005
R2886 VSS.n1995 VSS.n343 25.6005
R2887 VSS.n1995 VSS.n1994 25.6005
R2888 VSS.n1994 VSS.n345 25.6005
R2889 VSS.n1989 VSS.n345 25.6005
R2890 VSS.n1989 VSS.n1988 25.6005
R2891 VSS.n1988 VSS.n1987 25.6005
R2892 VSS.n1987 VSS.n347 25.6005
R2893 VSS.n1981 VSS.n347 25.6005
R2894 VSS.n1981 VSS.n1980 25.6005
R2895 VSS.n1980 VSS.n1979 25.6005
R2896 VSS.n1979 VSS.n349 25.6005
R2897 VSS.n1973 VSS.n349 25.6005
R2898 VSS.n1965 VSS.n1964 25.6005
R2899 VSS.n360 VSS.n357 25.6005
R2900 VSS.n1950 VSS.n1949 25.6005
R2901 VSS.n1949 VSS.n364 25.6005
R2902 VSS.n1944 VSS.n364 25.6005
R2903 VSS.n1944 VSS.n1943 25.6005
R2904 VSS.n1943 VSS.n1942 25.6005
R2905 VSS.n1942 VSS.n366 25.6005
R2906 VSS.n1936 VSS.n366 25.6005
R2907 VSS.n1936 VSS.n1935 25.6005
R2908 VSS.n1935 VSS.n1934 25.6005
R2909 VSS.n1934 VSS.n368 25.6005
R2910 VSS.n1928 VSS.n368 25.6005
R2911 VSS.n1928 VSS.n1927 25.6005
R2912 VSS.n1927 VSS.n1926 25.6005
R2913 VSS.n1926 VSS.n370 25.6005
R2914 VSS.n1920 VSS.n370 25.6005
R2915 VSS.n1836 VSS.n1834 25.6005
R2916 VSS.n1836 VSS.n1835 25.6005
R2917 VSS.n1835 VSS.n371 25.6005
R2918 VSS.n1848 VSS.n371 25.6005
R2919 VSS.n1849 VSS.n1848 25.6005
R2920 VSS.n1851 VSS.n1849 25.6005
R2921 VSS.n1852 VSS.n1851 25.6005
R2922 VSS.n1853 VSS.n1852 25.6005
R2923 VSS.n1854 VSS.n1853 25.6005
R2924 VSS.n1856 VSS.n1854 25.6005
R2925 VSS.n1857 VSS.n1856 25.6005
R2926 VSS.n1858 VSS.n1857 25.6005
R2927 VSS.n1859 VSS.n1858 25.6005
R2928 VSS.n1861 VSS.n1859 25.6005
R2929 VSS.n1862 VSS.n1861 25.6005
R2930 VSS.n1863 VSS.n1862 25.6005
R2931 VSS.n1864 VSS.n1863 25.6005
R2932 VSS.n1866 VSS.n1864 25.6005
R2933 VSS.n1867 VSS.n1866 25.6005
R2934 VSS.n1868 VSS.n1867 25.6005
R2935 VSS.n1869 VSS.n1868 25.6005
R2936 VSS.n1871 VSS.n1869 25.6005
R2937 VSS.n1872 VSS.n1871 25.6005
R2938 VSS.n1873 VSS.n1872 25.6005
R2939 VSS.n1874 VSS.n1873 25.6005
R2940 VSS.n1876 VSS.n1874 25.6005
R2941 VSS.n1877 VSS.n1876 25.6005
R2942 VSS.n1878 VSS.n1877 25.6005
R2943 VSS.n1879 VSS.n1878 25.6005
R2944 VSS.n1881 VSS.n1879 25.6005
R2945 VSS.n1882 VSS.n1881 25.6005
R2946 VSS.n1883 VSS.n1882 25.6005
R2947 VSS.n1884 VSS.n1883 25.6005
R2948 VSS.n1886 VSS.n1884 25.6005
R2949 VSS.n1887 VSS.n1886 25.6005
R2950 VSS.n1888 VSS.n1887 25.6005
R2951 VSS.n1889 VSS.n1888 25.6005
R2952 VSS.n1891 VSS.n1889 25.6005
R2953 VSS.n1892 VSS.n1891 25.6005
R2954 VSS.n1893 VSS.n1892 25.6005
R2955 VSS.n1894 VSS.n1893 25.6005
R2956 VSS.n1896 VSS.n1894 25.6005
R2957 VSS.n1897 VSS.n1896 25.6005
R2958 VSS.n1898 VSS.n1897 25.6005
R2959 VSS.n1899 VSS.n1898 25.6005
R2960 VSS.n1901 VSS.n1899 25.6005
R2961 VSS.n1902 VSS.n1901 25.6005
R2962 VSS.n1903 VSS.n1902 25.6005
R2963 VSS.n1904 VSS.n1903 25.6005
R2964 VSS.n1906 VSS.n1904 25.6005
R2965 VSS.n1907 VSS.n1906 25.6005
R2966 VSS.n1908 VSS.n1907 25.6005
R2967 VSS.n1909 VSS.n1908 25.6005
R2968 VSS.n1911 VSS.n1909 25.6005
R2969 VSS.n1912 VSS.n1911 25.6005
R2970 VSS.n1913 VSS.n1912 25.6005
R2971 VSS.n1914 VSS.n1913 25.6005
R2972 VSS.n1916 VSS.n1914 25.6005
R2973 VSS.n1917 VSS.n1916 25.6005
R2974 VSS.n1918 VSS.n1917 25.6005
R2975 VSS.n1919 VSS.n1918 25.6005
R2976 VSS.n1828 VSS.n1827 25.6005
R2977 VSS.n1827 VSS.n1826 25.6005
R2978 VSS.n1826 VSS.n1823 25.6005
R2979 VSS.n1823 VSS.n1822 25.6005
R2980 VSS.n1822 VSS.n1819 25.6005
R2981 VSS.n1819 VSS.n1818 25.6005
R2982 VSS.n1818 VSS.n1815 25.6005
R2983 VSS.n1815 VSS.n1814 25.6005
R2984 VSS.n1814 VSS.n1811 25.6005
R2985 VSS.n1811 VSS.n1810 25.6005
R2986 VSS.n1810 VSS.n1807 25.6005
R2987 VSS.n1807 VSS.n1806 25.6005
R2988 VSS.n1806 VSS.n1803 25.6005
R2989 VSS.n1803 VSS.n1802 25.6005
R2990 VSS.n1794 VSS.n1791 25.6005
R2991 VSS.n407 VSS.n403 25.6005
R2992 VSS.n1780 VSS.n1779 25.6005
R2993 VSS.n1779 VSS.n1776 25.6005
R2994 VSS.n1776 VSS.n1775 25.6005
R2995 VSS.n1775 VSS.n1772 25.6005
R2996 VSS.n1772 VSS.n1771 25.6005
R2997 VSS.n1771 VSS.n1768 25.6005
R2998 VSS.n1768 VSS.n1767 25.6005
R2999 VSS.n1767 VSS.n1764 25.6005
R3000 VSS.n1764 VSS.n1763 25.6005
R3001 VSS.n1763 VSS.n1760 25.6005
R3002 VSS.n1760 VSS.n1759 25.6005
R3003 VSS.n1759 VSS.n1756 25.6005
R3004 VSS.n1756 VSS.n1755 25.6005
R3005 VSS.n1755 VSS.n378 25.6005
R3006 VSS.n1833 VSS.n378 25.6005
R3007 VSS.n945 VSS.n574 25.6005
R3008 VSS.n945 VSS.n944 25.6005
R3009 VSS.n951 VSS.n944 25.6005
R3010 VSS.n952 VSS.n951 25.6005
R3011 VSS.n953 VSS.n952 25.6005
R3012 VSS.n953 VSS.n942 25.6005
R3013 VSS.n959 VSS.n942 25.6005
R3014 VSS.n960 VSS.n959 25.6005
R3015 VSS.n961 VSS.n960 25.6005
R3016 VSS.n961 VSS.n940 25.6005
R3017 VSS.n967 VSS.n940 25.6005
R3018 VSS.n968 VSS.n967 25.6005
R3019 VSS.n969 VSS.n968 25.6005
R3020 VSS.n969 VSS.n938 25.6005
R3021 VSS.n975 VSS.n938 25.6005
R3022 VSS.n976 VSS.n975 25.6005
R3023 VSS.n977 VSS.n976 25.6005
R3024 VSS.n977 VSS.n936 25.6005
R3025 VSS.n982 VSS.n936 25.6005
R3026 VSS.n983 VSS.n982 25.6005
R3027 VSS.n983 VSS.n934 25.6005
R3028 VSS.n988 VSS.n934 25.6005
R3029 VSS.n1626 VSS.n1625 25.6005
R3030 VSS.n1625 VSS.n1624 25.6005
R3031 VSS.n1624 VSS.n575 25.6005
R3032 VSS.n590 VSS.n575 25.6005
R3033 VSS.n1612 VSS.n590 25.6005
R3034 VSS.n1612 VSS.n1611 25.6005
R3035 VSS.n1611 VSS.n1610 25.6005
R3036 VSS.n1610 VSS.n591 25.6005
R3037 VSS.n605 VSS.n591 25.6005
R3038 VSS.n1598 VSS.n605 25.6005
R3039 VSS.n1598 VSS.n1597 25.6005
R3040 VSS.n1596 VSS.n606 25.6005
R3041 VSS.n1591 VSS.n606 25.6005
R3042 VSS.n1591 VSS.n1590 25.6005
R3043 VSS.n1590 VSS.n1589 25.6005
R3044 VSS.n1589 VSS.n1586 25.6005
R3045 VSS.n1586 VSS.n1585 25.6005
R3046 VSS.n1585 VSS.n1582 25.6005
R3047 VSS.n1582 VSS.n1581 25.6005
R3048 VSS.n1581 VSS.n1578 25.6005
R3049 VSS.n1578 VSS.n1577 25.6005
R3050 VSS.n1577 VSS.n1574 25.6005
R3051 VSS.n1574 VSS.n1573 25.6005
R3052 VSS.n1573 VSS.n1570 25.6005
R3053 VSS.n1570 VSS.n1569 25.6005
R3054 VSS.n1569 VSS.n1566 25.6005
R3055 VSS.n1566 VSS.n1565 25.6005
R3056 VSS.n1565 VSS.n1562 25.6005
R3057 VSS.n1562 VSS.n1561 25.6005
R3058 VSS.n1561 VSS.n1558 25.6005
R3059 VSS.n1558 VSS.n1557 25.6005
R3060 VSS.n1557 VSS.n1554 25.6005
R3061 VSS.n1554 VSS.n1553 25.6005
R3062 VSS.n1066 VSS.n989 25.6005
R3063 VSS.n1062 VSS.n1059 25.6005
R3064 VSS.n997 VSS.n995 25.6005
R3065 VSS.n1000 VSS.n999 25.6005
R3066 VSS.n999 VSS.n620 25.6005
R3067 VSS.n1342 VSS.n715 25.6005
R3068 VSS.n1359 VSS.n715 25.6005
R3069 VSS.n1360 VSS.n1359 25.6005
R3070 VSS.n1361 VSS.n1360 25.6005
R3071 VSS.n1361 VSS.n705 25.6005
R3072 VSS.n1416 VSS.n705 25.6005
R3073 VSS.n1416 VSS.n1415 25.6005
R3074 VSS.n1415 VSS.n1414 25.6005
R3075 VSS.n1414 VSS.n706 25.6005
R3076 VSS.n706 VSS.n510 25.6005
R3077 VSS.n1642 VSS.n510 25.6005
R3078 VSS.n1341 VSS.n1340 25.6005
R3079 VSS.n1340 VSS.n1280 25.6005
R3080 VSS.n1281 VSS.n1280 25.6005
R3081 VSS.n1333 VSS.n1281 25.6005
R3082 VSS.n1333 VSS.n1332 25.6005
R3083 VSS.n1332 VSS.n1331 25.6005
R3084 VSS.n1331 VSS.n1283 25.6005
R3085 VSS.n1326 VSS.n1283 25.6005
R3086 VSS.n1326 VSS.n1325 25.6005
R3087 VSS.n1325 VSS.n1324 25.6005
R3088 VSS.n1324 VSS.n1286 25.6005
R3089 VSS.n1319 VSS.n1286 25.6005
R3090 VSS.n1319 VSS.n1318 25.6005
R3091 VSS.n1318 VSS.n1317 25.6005
R3092 VSS.n1317 VSS.n1289 25.6005
R3093 VSS.n1312 VSS.n1289 25.6005
R3094 VSS.n1312 VSS.n1311 25.6005
R3095 VSS.n1311 VSS.n1310 25.6005
R3096 VSS.n1310 VSS.n1292 25.6005
R3097 VSS.n1305 VSS.n1292 25.6005
R3098 VSS.n1305 VSS.n1304 25.6005
R3099 VSS.n1304 VSS.n1303 25.6005
R3100 VSS.n1300 VSS.n1299 25.6005
R3101 VSS.n1299 VSS.n1297 25.6005
R3102 VSS.n1297 VSS.n1296 25.6005
R3103 VSS.n1296 VSS.n711 25.6005
R3104 VSS.n1367 VSS.n711 25.6005
R3105 VSS.n1368 VSS.n1367 25.6005
R3106 VSS.n1374 VSS.n504 25.6005
R3107 VSS.n1641 VSS.n1640 25.6005
R3108 VSS.n1640 VSS.n511 25.6005
R3109 VSS.n525 VSS.n511 25.6005
R3110 VSS.n526 VSS.n525 25.6005
R3111 VSS.n529 VSS.n526 25.6005
R3112 VSS.n530 VSS.n529 25.6005
R3113 VSS.n533 VSS.n530 25.6005
R3114 VSS.n534 VSS.n533 25.6005
R3115 VSS.n537 VSS.n534 25.6005
R3116 VSS.n538 VSS.n537 25.6005
R3117 VSS.n541 VSS.n538 25.6005
R3118 VSS.n542 VSS.n541 25.6005
R3119 VSS.n545 VSS.n542 25.6005
R3120 VSS.n546 VSS.n545 25.6005
R3121 VSS.n549 VSS.n546 25.6005
R3122 VSS.n550 VSS.n549 25.6005
R3123 VSS.n553 VSS.n550 25.6005
R3124 VSS.n554 VSS.n553 25.6005
R3125 VSS.n557 VSS.n554 25.6005
R3126 VSS.n558 VSS.n557 25.6005
R3127 VSS.n560 VSS.n558 25.6005
R3128 VSS.n560 VSS.n559 25.6005
R3129 VSS.n2143 VSS.n2142 25.6005
R3130 VSS.n2142 VSS.n2135 25.6005
R3131 VSS.n2136 VSS.n2135 25.6005
R3132 VSS.n2136 VSS.n2131 25.6005
R3133 VSS.n2144 VSS.n2127 25.6005
R3134 VSS.n2154 VSS.n2127 25.6005
R3135 VSS.n2155 VSS.n2154 25.6005
R3136 VSS.n2156 VSS.n2155 25.6005
R3137 VSS.n2156 VSS.n2119 25.6005
R3138 VSS.n2167 VSS.n2119 25.6005
R3139 VSS.n2168 VSS.n2167 25.6005
R3140 VSS.n2169 VSS.n2168 25.6005
R3141 VSS.n2169 VSS.n233 25.6005
R3142 VSS.n2179 VSS.n233 25.6005
R3143 VSS.n2180 VSS.n2179 25.6005
R3144 VSS.n2181 VSS.n2180 25.6005
R3145 VSS.n2181 VSS.n225 25.6005
R3146 VSS.n2191 VSS.n225 25.6005
R3147 VSS.n2192 VSS.n2191 25.6005
R3148 VSS.n2193 VSS.n2192 25.6005
R3149 VSS.n2193 VSS.n217 25.6005
R3150 VSS.n2203 VSS.n217 25.6005
R3151 VSS.n2204 VSS.n2203 25.6005
R3152 VSS.n2205 VSS.n2204 25.6005
R3153 VSS.n2205 VSS.n209 25.6005
R3154 VSS.n2215 VSS.n209 25.6005
R3155 VSS.n2216 VSS.n2215 25.6005
R3156 VSS.n2217 VSS.n2216 25.6005
R3157 VSS.n2217 VSS.n201 25.6005
R3158 VSS.n2227 VSS.n201 25.6005
R3159 VSS.n2228 VSS.n2227 25.6005
R3160 VSS.n2229 VSS.n2228 25.6005
R3161 VSS.n2229 VSS.n192 25.6005
R3162 VSS.n2239 VSS.n192 25.6005
R3163 VSS.n2240 VSS.n2239 25.6005
R3164 VSS.n2241 VSS.n2240 25.6005
R3165 VSS.n2241 VSS.n184 25.6005
R3166 VSS.n2251 VSS.n184 25.6005
R3167 VSS.n2252 VSS.n2251 25.6005
R3168 VSS.n2253 VSS.n2252 25.6005
R3169 VSS.n2253 VSS.n176 25.6005
R3170 VSS.n2263 VSS.n176 25.6005
R3171 VSS.n2264 VSS.n2263 25.6005
R3172 VSS.n2265 VSS.n2264 25.6005
R3173 VSS.n2265 VSS.n168 25.6005
R3174 VSS.n2275 VSS.n168 25.6005
R3175 VSS.n2276 VSS.n2275 25.6005
R3176 VSS.n2277 VSS.n2276 25.6005
R3177 VSS.n2277 VSS.n160 25.6005
R3178 VSS.n2287 VSS.n160 25.6005
R3179 VSS.n2288 VSS.n2287 25.6005
R3180 VSS.n2289 VSS.n2288 25.6005
R3181 VSS.n2289 VSS.n152 25.6005
R3182 VSS.n2300 VSS.n152 25.6005
R3183 VSS.n2301 VSS.n2300 25.6005
R3184 VSS.n2302 VSS.n2301 25.6005
R3185 VSS.n2302 VSS.n138 25.6005
R3186 VSS.n2310 VSS.n146 25.6005
R3187 VSS.n2310 VSS.n2309 25.6005
R3188 VSS.n2309 VSS.n2308 25.6005
R3189 VSS.n2149 VSS.n2148 25.6005
R3190 VSS.n2150 VSS.n2149 25.6005
R3191 VSS.n2150 VSS.n2123 25.6005
R3192 VSS.n2160 VSS.n2123 25.6005
R3193 VSS.n2161 VSS.n2160 25.6005
R3194 VSS.n2162 VSS.n2161 25.6005
R3195 VSS.n2162 VSS.n237 25.6005
R3196 VSS.n2173 VSS.n237 25.6005
R3197 VSS.n2174 VSS.n2173 25.6005
R3198 VSS.n2175 VSS.n2174 25.6005
R3199 VSS.n2175 VSS.n229 25.6005
R3200 VSS.n2185 VSS.n229 25.6005
R3201 VSS.n2186 VSS.n2185 25.6005
R3202 VSS.n2187 VSS.n2186 25.6005
R3203 VSS.n2187 VSS.n221 25.6005
R3204 VSS.n2197 VSS.n221 25.6005
R3205 VSS.n2198 VSS.n2197 25.6005
R3206 VSS.n2199 VSS.n2198 25.6005
R3207 VSS.n2199 VSS.n213 25.6005
R3208 VSS.n2209 VSS.n213 25.6005
R3209 VSS.n2210 VSS.n2209 25.6005
R3210 VSS.n2211 VSS.n2210 25.6005
R3211 VSS.n2211 VSS.n205 25.6005
R3212 VSS.n2221 VSS.n205 25.6005
R3213 VSS.n2222 VSS.n2221 25.6005
R3214 VSS.n2223 VSS.n2222 25.6005
R3215 VSS.n2223 VSS.n196 25.6005
R3216 VSS.n2233 VSS.n196 25.6005
R3217 VSS.n2234 VSS.n2233 25.6005
R3218 VSS.n2235 VSS.n2234 25.6005
R3219 VSS.n2235 VSS.n188 25.6005
R3220 VSS.n2245 VSS.n188 25.6005
R3221 VSS.n2246 VSS.n2245 25.6005
R3222 VSS.n2247 VSS.n2246 25.6005
R3223 VSS.n2247 VSS.n180 25.6005
R3224 VSS.n2257 VSS.n180 25.6005
R3225 VSS.n2258 VSS.n2257 25.6005
R3226 VSS.n2259 VSS.n2258 25.6005
R3227 VSS.n2259 VSS.n172 25.6005
R3228 VSS.n2269 VSS.n172 25.6005
R3229 VSS.n2270 VSS.n2269 25.6005
R3230 VSS.n2271 VSS.n2270 25.6005
R3231 VSS.n2271 VSS.n164 25.6005
R3232 VSS.n2281 VSS.n164 25.6005
R3233 VSS.n2282 VSS.n2281 25.6005
R3234 VSS.n2283 VSS.n2282 25.6005
R3235 VSS.n2283 VSS.n156 25.6005
R3236 VSS.n2293 VSS.n156 25.6005
R3237 VSS.n2294 VSS.n2293 25.6005
R3238 VSS.n2296 VSS.n2294 25.6005
R3239 VSS.n2296 VSS.n2295 25.6005
R3240 VSS.n2295 VSS.n149 25.6005
R3241 VSS.n149 VSS.n147 25.6005
R3242 VSS.n1095 VSS.n1094 25.6005
R3243 VSS.n1096 VSS.n1095 25.6005
R3244 VSS.n1096 VSS.n768 25.6005
R3245 VSS.n1102 VSS.n768 25.6005
R3246 VSS.n1103 VSS.n1102 25.6005
R3247 VSS.n1104 VSS.n1103 25.6005
R3248 VSS.n1104 VSS.n766 25.6005
R3249 VSS.n1110 VSS.n766 25.6005
R3250 VSS.n1111 VSS.n1110 25.6005
R3251 VSS.n1112 VSS.n1111 25.6005
R3252 VSS.n1112 VSS.n764 25.6005
R3253 VSS.n1118 VSS.n764 25.6005
R3254 VSS.n1119 VSS.n1118 25.6005
R3255 VSS.n1120 VSS.n1119 25.6005
R3256 VSS.n1120 VSS.n762 25.6005
R3257 VSS.n1126 VSS.n762 25.6005
R3258 VSS.n1127 VSS.n1126 25.6005
R3259 VSS.n1128 VSS.n1127 25.6005
R3260 VSS.n1128 VSS.n760 25.6005
R3261 VSS.n1133 VSS.n760 25.6005
R3262 VSS.n1134 VSS.n1133 25.6005
R3263 VSS.n1137 VSS.n1134 25.6005
R3264 VSS.n1141 VSS.n1138 25.6005
R3265 VSS.n1142 VSS.n1141 25.6005
R3266 VSS.n1145 VSS.n1142 25.6005
R3267 VSS.n1146 VSS.n1145 25.6005
R3268 VSS.n1149 VSS.n1146 25.6005
R3269 VSS.n1150 VSS.n1149 25.6005
R3270 VSS.n1153 VSS.n1150 25.6005
R3271 VSS.n1154 VSS.n1153 25.6005
R3272 VSS.n1157 VSS.n1154 25.6005
R3273 VSS.n1158 VSS.n1157 25.6005
R3274 VSS.n1161 VSS.n1158 25.6005
R3275 VSS.n1162 VSS.n1161 25.6005
R3276 VSS.n1165 VSS.n1162 25.6005
R3277 VSS.n1166 VSS.n1165 25.6005
R3278 VSS.n1169 VSS.n1166 25.6005
R3279 VSS.n1170 VSS.n1169 25.6005
R3280 VSS.n1173 VSS.n1170 25.6005
R3281 VSS.n1174 VSS.n1173 25.6005
R3282 VSS.n1177 VSS.n1174 25.6005
R3283 VSS.n1178 VSS.n1177 25.6005
R3284 VSS.n1181 VSS.n1178 25.6005
R3285 VSS.n1182 VSS.n1181 25.6005
R3286 VSS.n1185 VSS.n1182 25.6005
R3287 VSS.n1189 VSS.n1186 25.6005
R3288 VSS.n1190 VSS.n1189 25.6005
R3289 VSS.n1193 VSS.n1190 25.6005
R3290 VSS.n1194 VSS.n1193 25.6005
R3291 VSS.n1197 VSS.n1194 25.6005
R3292 VSS.n1198 VSS.n1197 25.6005
R3293 VSS.n1201 VSS.n1198 25.6005
R3294 VSS.n1202 VSS.n1201 25.6005
R3295 VSS.n1205 VSS.n1202 25.6005
R3296 VSS.n1206 VSS.n1205 25.6005
R3297 VSS.n1209 VSS.n1206 25.6005
R3298 VSS.n1210 VSS.n1209 25.6005
R3299 VSS.n1213 VSS.n1210 25.6005
R3300 VSS.n1214 VSS.n1213 25.6005
R3301 VSS.n1217 VSS.n1214 25.6005
R3302 VSS.n1218 VSS.n1217 25.6005
R3303 VSS.n1221 VSS.n1218 25.6005
R3304 VSS.n1222 VSS.n1221 25.6005
R3305 VSS.n1225 VSS.n1222 25.6005
R3306 VSS.n1226 VSS.n1225 25.6005
R3307 VSS.n1229 VSS.n1226 25.6005
R3308 VSS.n1230 VSS.n1229 25.6005
R3309 VSS.n1233 VSS.n1230 25.6005
R3310 VSS.n1237 VSS.n1234 25.6005
R3311 VSS.n1238 VSS.n1237 25.6005
R3312 VSS.n1241 VSS.n1238 25.6005
R3313 VSS.n1242 VSS.n1241 25.6005
R3314 VSS.n1245 VSS.n1242 25.6005
R3315 VSS.n1246 VSS.n1245 25.6005
R3316 VSS.n1249 VSS.n1246 25.6005
R3317 VSS.n1250 VSS.n1249 25.6005
R3318 VSS.n1253 VSS.n1250 25.6005
R3319 VSS.n1254 VSS.n1253 25.6005
R3320 VSS.n1257 VSS.n1254 25.6005
R3321 VSS.n1258 VSS.n1257 25.6005
R3322 VSS.n1261 VSS.n1258 25.6005
R3323 VSS.n1262 VSS.n1261 25.6005
R3324 VSS.n1265 VSS.n1262 25.6005
R3325 VSS.n1266 VSS.n1265 25.6005
R3326 VSS.n1269 VSS.n1266 25.6005
R3327 VSS.n1271 VSS.n1269 25.6005
R3328 VSS.n1272 VSS.n1271 25.6005
R3329 VSS.n1273 VSS.n1272 25.6005
R3330 VSS.n1273 VSS.n721 25.6005
R3331 VSS.n1348 VSS.n721 25.6005
R3332 VSS.n1086 VSS.n1085 25.6005
R3333 VSS.n906 VSS.n775 25.6005
R3334 VSS.n910 VSS.n898 25.6005
R3335 VSS.n899 VSS.n894 25.6005
R3336 VSS.n918 VSS.n894 25.6005
R3337 VSS.n919 VSS.n918 25.6005
R3338 VSS.n920 VSS.n919 25.6005
R3339 VSS.n920 VSS.n890 25.6005
R3340 VSS.n926 VSS.n890 25.6005
R3341 VSS.n927 VSS.n926 25.6005
R3342 VSS.n929 VSS.n882 25.6005
R3343 VSS.n1075 VSS.n882 25.6005
R3344 VSS.n1075 VSS.n883 25.6005
R3345 VSS.n1016 VSS.n883 25.6005
R3346 VSS.n1018 VSS.n1006 25.6005
R3347 VSS.n1046 VSS.n1006 25.6005
R3348 VSS.n1046 VSS.n1045 25.6005
R3349 VSS.n1045 VSS.n1044 25.6005
R3350 VSS.n1044 VSS.n1007 25.6005
R3351 VSS.n1009 VSS.n1007 25.6005
R3352 VSS.n1012 VSS.n1009 25.6005
R3353 VSS.n1034 VSS.n1033 25.6005
R3354 VSS.n2351 VSS.n125 25.6005
R3355 VSS.n2357 VSS.n119 25.6005
R3356 VSS.n2395 VSS.n2394 25.6005
R3357 VSS.n2394 VSS.n2393 25.6005
R3358 VSS.n2393 VSS.n2392 25.6005
R3359 VSS.n2392 VSS.n2390 25.6005
R3360 VSS.n2390 VSS.n2387 25.6005
R3361 VSS.n2387 VSS.n2386 25.6005
R3362 VSS.n2386 VSS.n2383 25.6005
R3363 VSS.n2383 VSS.n2382 25.6005
R3364 VSS.n2382 VSS.n2379 25.6005
R3365 VSS.n2379 VSS.n2378 25.6005
R3366 VSS.n2378 VSS.n2375 25.6005
R3367 VSS.n2375 VSS.n2374 25.6005
R3368 VSS.n2374 VSS.n2371 25.6005
R3369 VSS.n2371 VSS.n2370 25.6005
R3370 VSS.n2370 VSS.n2367 25.6005
R3371 VSS.n2367 VSS.n2366 25.6005
R3372 VSS.n2366 VSS.n2363 25.6005
R3373 VSS.n2363 VSS.n2362 25.6005
R3374 VSS.n2362 VSS.n104 25.6005
R3375 VSS.n104 VSS.n102 25.6005
R3376 VSS.n2403 VSS.n102 25.6005
R3377 VSS.n2404 VSS.n2403 25.6005
R3378 VSS.n2405 VSS.n100 25.6005
R3379 VSS.n2411 VSS.n100 25.6005
R3380 VSS.n2412 VSS.n2411 25.6005
R3381 VSS.n2413 VSS.n2412 25.6005
R3382 VSS.n2413 VSS.n98 25.6005
R3383 VSS.n2419 VSS.n98 25.6005
R3384 VSS.n2420 VSS.n2419 25.6005
R3385 VSS.n2421 VSS.n2420 25.6005
R3386 VSS.n2421 VSS.n96 25.6005
R3387 VSS.n2427 VSS.n96 25.6005
R3388 VSS.n2428 VSS.n2427 25.6005
R3389 VSS.n2429 VSS.n2428 25.6005
R3390 VSS.n2429 VSS.n94 25.6005
R3391 VSS.n2435 VSS.n94 25.6005
R3392 VSS.n2436 VSS.n2435 25.6005
R3393 VSS.n2437 VSS.n2436 25.6005
R3394 VSS.n2437 VSS.n92 25.6005
R3395 VSS.n2443 VSS.n92 25.6005
R3396 VSS.n2444 VSS.n2443 25.6005
R3397 VSS.n2445 VSS.n2444 25.6005
R3398 VSS.n2445 VSS.n90 25.6005
R3399 VSS.n2451 VSS.n90 25.6005
R3400 VSS.n2452 VSS.n2451 25.6005
R3401 VSS.n2453 VSS.n88 25.6005
R3402 VSS.n2459 VSS.n88 25.6005
R3403 VSS.n2460 VSS.n2459 25.6005
R3404 VSS.n2461 VSS.n2460 25.6005
R3405 VSS.n2461 VSS.n86 25.6005
R3406 VSS.n2467 VSS.n86 25.6005
R3407 VSS.n2468 VSS.n2467 25.6005
R3408 VSS.n2469 VSS.n2468 25.6005
R3409 VSS.n2469 VSS.n84 25.6005
R3410 VSS.n2475 VSS.n84 25.6005
R3411 VSS.n2476 VSS.n2475 25.6005
R3412 VSS.n2477 VSS.n2476 25.6005
R3413 VSS.n2477 VSS.n82 25.6005
R3414 VSS.n2483 VSS.n82 25.6005
R3415 VSS.n2484 VSS.n2483 25.6005
R3416 VSS.n2485 VSS.n2484 25.6005
R3417 VSS.n2485 VSS.n80 25.6005
R3418 VSS.n2491 VSS.n80 25.6005
R3419 VSS.n2492 VSS.n2491 25.6005
R3420 VSS.n2493 VSS.n2492 25.6005
R3421 VSS.n2493 VSS.n78 25.6005
R3422 VSS.n2499 VSS.n78 25.6005
R3423 VSS.n2500 VSS.n2499 25.6005
R3424 VSS.n2501 VSS.n76 25.6005
R3425 VSS.n2507 VSS.n76 25.6005
R3426 VSS.n2508 VSS.n2507 25.6005
R3427 VSS.n2509 VSS.n2508 25.6005
R3428 VSS.n2509 VSS.n74 25.6005
R3429 VSS.n2515 VSS.n74 25.6005
R3430 VSS.n2516 VSS.n2515 25.6005
R3431 VSS.n2517 VSS.n2516 25.6005
R3432 VSS.n2517 VSS.n72 25.6005
R3433 VSS.n2523 VSS.n72 25.6005
R3434 VSS.n2524 VSS.n2523 25.6005
R3435 VSS.n2525 VSS.n2524 25.6005
R3436 VSS.n2525 VSS.n70 25.6005
R3437 VSS.n2531 VSS.n70 25.6005
R3438 VSS.n2532 VSS.n2531 25.6005
R3439 VSS.n2533 VSS.n2532 25.6005
R3440 VSS.n2533 VSS.n68 25.6005
R3441 VSS.n2539 VSS.n68 25.6005
R3442 VSS.n2540 VSS.n2539 25.6005
R3443 VSS.n2541 VSS.n2540 25.6005
R3444 VSS.n2541 VSS.n66 25.6005
R3445 VSS.n66 VSS.n64 25.6005
R3446 VSS.n1351 VSS.n697 25.6005
R3447 VSS.n1421 VSS.n698 25.6005
R3448 VSS.n1409 VSS.n1381 25.6005
R3449 VSS.n1387 VSS.n1386 25.6005
R3450 VSS.n1386 VSS.n1382 25.6005
R3451 VSS.n1382 VSS.n566 25.6005
R3452 VSS.n1634 VSS.n566 25.6005
R3453 VSS.n1634 VSS.n1633 25.6005
R3454 VSS.n1633 VSS.n1632 25.6005
R3455 VSS.n1632 VSS.n567 25.6005
R3456 VSS.n1619 VSS.n581 25.6005
R3457 VSS.n1619 VSS.n1618 25.6005
R3458 VSS.n1618 VSS.n1617 25.6005
R3459 VSS.n1617 VSS.n583 25.6005
R3460 VSS.n1605 VSS.n1604 25.6005
R3461 VSS.n1604 VSS.n1603 25.6005
R3462 VSS.n1603 VSS.n599 25.6005
R3463 VSS.n1547 VSS.n599 25.6005
R3464 VSS.n1547 VSS.n1546 25.6005
R3465 VSS.n1546 VSS.n1545 25.6005
R3466 VSS.n1545 VSS.n622 25.6005
R3467 VSS.n649 VSS.n647 25.6005
R3468 VSS.n1491 VSS.n1490 25.6005
R3469 VSS.n2554 VSS.n2553 25.6005
R3470 VSS.n2599 VSS.t59 25.0064
R3471 VSS.n2171 VSS.n2117 24.8841
R3472 VSS.n687 VSS.n657 24.8476
R3473 VSS.n1445 VSS.n1443 24.8476
R3474 VSS.n827 VSS.n826 24.8476
R3475 VSS.n853 VSS.n850 24.8476
R3476 VSS.n471 VSS.n453 24.8476
R3477 VSS.n425 VSS.n424 24.8476
R3478 VSS.n1669 VSS.n1663 24.8476
R3479 VSS.n1724 VSS.n1718 24.8476
R3480 VSS.n1957 VSS.n1956 24.8476
R3481 VSS.n1784 VSS.n1783 24.8476
R3482 VSS.n1647 VSS.n1646 24.8476
R3483 VSS.n931 VSS.n930 24.8476
R3484 VSS.n1025 VSS.n1024 24.8476
R3485 VSS.n1399 VSS.n1398 24.8476
R3486 VSS.n1390 VSS.n1389 24.8476
R3487 VSS.n466 VSS.n465 24.75
R3488 VSS.n429 VSS.n428 24.75
R3489 VSS.n459 VSS.n455 24.2609
R3490 VSS.n433 VSS.n412 24.2609
R3491 VSS.n1682 VSS.n1658 24.2609
R3492 VSS.n1676 VSS.n1656 24.2609
R3493 VSS.n1737 VSS.n1731 24.2609
R3494 VSS.n1742 VSS.n1733 24.2609
R3495 VSS.n1972 VSS.n351 23.7181
R3496 VSS.n1969 VSS.n353 23.7181
R3497 VSS.n1799 VSS.n399 23.7181
R3498 VSS.n1795 VSS.n400 23.7181
R3499 VSS.n2316 VSS.n2315 23.7181
R3500 VSS.n1637 VSS.n1636 23.4436
R3501 VSS.n686 VSS.n659 23.3417
R3502 VSS.n1449 VSS.n1448 23.3417
R3503 VSS.n823 VSS.n797 23.3417
R3504 VSS.n854 VSS.n848 23.3417
R3505 VSS.n475 VSS.n474 23.3417
R3506 VSS.n459 VSS.n456 23.3417
R3507 VSS.n434 VSS.n433 23.3417
R3508 VSS.n421 VSS.n416 23.3417
R3509 VSS.n1682 VSS.n1659 23.3417
R3510 VSS.n1676 VSS.n1657 23.3417
R3511 VSS.n1666 VSS.n1662 23.3417
R3512 VSS.n1737 VSS.n1732 23.3417
R3513 VSS.n1742 VSS.n1734 23.3417
R3514 VSS.n1721 VSS.n1717 23.3417
R3515 VSS.n2609 VSS.n2603 22.9652
R3516 VSS.n909 VSS.n899 22.9652
R3517 VSS.n1013 VSS.n1012 22.9652
R3518 VSS.n1408 VSS.n1387 22.9652
R3519 VSS.n650 VSS.n622 22.9652
R3520 VSS.n1493 VSS.n644 22.9226
R3521 VSS.n2556 VSS.n57 22.9226
R3522 VSS.n2546 VSS.n52 22.9226
R3523 VSS.n1670 VSS.n1669 22.4252
R3524 VSS.n1725 VSS.n1724 22.4252
R3525 VSS.n2108 VSS.t5 22.4016
R3526 VSS.t0 VSS.n2021 22.4016
R3527 VSS.n683 VSS.n682 21.8358
R3528 VSS.n1452 VSS.n1441 21.8358
R3529 VSS.n822 VSS.n799 21.8358
R3530 VSS.n858 VSS.n857 21.8358
R3531 VSS.n477 VSS.n451 21.8358
R3532 VSS.n463 VSS.n462 21.8358
R3533 VSS.n436 VSS.n411 21.8358
R3534 VSS.n420 VSS.n417 21.8358
R3535 VSS.n1686 VSS.n1685 21.8358
R3536 VSS.n1689 VSS.n1655 21.8358
R3537 VSS.n1672 VSS.n1661 21.8358
R3538 VSS.n1749 VSS.n1730 21.8358
R3539 VSS.n1746 VSS.n1745 21.8358
R3540 VSS.n1727 VSS.n1716 21.8358
R3541 VSS.n1065 VSS.n990 21.8358
R3542 VSS.n1373 VSS.n1372 21.8358
R3543 VSS.n907 VSS.n906 21.8358
R3544 VSS.n1032 VSS.n125 21.8358
R3545 VSS.n1406 VSS.n698 21.8358
R3546 VSS.n1491 VSS.n1489 21.8358
R3547 VSS.n2069 VSS.t14 21.3597
R3548 VSS.t26 VSS.n2060 21.3597
R3549 VSS.n1961 VSS.n355 21.0829
R3550 VSS.n1956 VSS.n361 21.0829
R3551 VSS.n1788 VSS.n402 21.0829
R3552 VSS.n1783 VSS.n408 21.0829
R3553 VSS.n1085 VSS.n1084 21.0829
R3554 VSS.n2350 VSS.n119 21.0829
R3555 VSS.n1422 VSS.n697 21.0829
R3556 VSS.n2554 VSS.n61 21.0829
R3557 VSS.n1069 VSS.n886 20.4928
R3558 VSS.n679 VSS.n661 20.3299
R3559 VSS.n1453 VSS.n1439 20.3299
R3560 VSS.n819 VSS.n818 20.3299
R3561 VSS.n861 VSS.n846 20.3299
R3562 VSS.n777 VSS.n774 20.3299
R3563 VSS.n2358 VSS.n117 20.3299
R3564 VSS.n1354 VSS.n1353 20.3299
R3565 VSS.n2552 VSS.n62 20.3299
R3566 VSS.n260 VSS.t34 20.3178
R3567 VSS.n2030 VSS.t38 20.3178
R3568 VSS.n2563 VSS.t2 20.3178
R3569 VSS.n1961 VSS.n1960 19.9534
R3570 VSS.n1788 VSS.n1787 19.9534
R3571 VSS.n1629 VSS.n1628 19.7969
R3572 VSS.n1068 VSS.n571 19.7969
R3573 VSS.n1621 VSS.n578 19.7969
R3574 VSS.n586 VSS.n585 19.7969
R3575 VSS.n1615 VSS.n1614 19.7969
R3576 VSS.n1608 VSS.n593 19.7969
R3577 VSS.n1607 VSS.n595 19.7969
R3578 VSS.n1049 VSS.n1001 19.7969
R3579 VSS.n1601 VSS.n1600 19.7969
R3580 VSS.n1550 VSS.n602 19.7969
R3581 VSS.n678 VSS.n663 18.824
R3582 VSS.n1457 VSS.n1456 18.824
R3583 VSS.n815 VSS.n801 18.824
R3584 VSS.n862 VSS.n844 18.824
R3585 VSS.n1371 VSS.n710 18.824
R3586 VSS.n1278 VSS.n1277 18.7549
R3587 VSS.n1357 VSS.n1356 18.7549
R3588 VSS.n1364 VSS.n1363 18.7549
R3589 VSS.n1418 VSS.n702 18.7549
R3590 VSS.n1412 VSS.n1411 18.7549
R3591 VSS.n1378 VSS.n507 18.7549
R3592 VSS.n1646 VSS.n503 18.5363
R3593 VSS.n2608 VSS.n2607 18.4476
R3594 VSS.n928 VSS.n927 18.4476
R3595 VSS.n1018 VSS.n1015 18.4476
R3596 VSS.n1396 VSS.n567 18.4476
R3597 VSS.n1605 VSS.n598 18.4476
R3598 VSS.n1543 VSS.t10 18.234
R3599 VSS.n26 VSS.n16 18.0711
R3600 VSS.n1052 VSS.n998 18.0711
R3601 VSS.n1365 VSS.t18 17.713
R3602 VSS.n993 VSS.t12 17.713
R3603 VSS.n2569 VSS.t19 17.713
R3604 VSS.n675 VSS.n674 17.3181
R3605 VSS.n1460 VSS.n1437 17.3181
R3606 VSS.n814 VSS.n803 17.3181
R3607 VSS.n867 VSS.n866 17.3181
R3608 VSS.n1970 VSS.n1969 17.3181
R3609 VSS.n1798 VSS.n400 17.3181
R3610 VSS.n1063 VSS.n1062 17.3181
R3611 VSS.n668 VSS.n667 17.1928
R3612 VSS.n1465 VSS.n1433 17.1928
R3613 VSS.n807 VSS.n806 17.1928
R3614 VSS.n873 VSS.n872 17.1928
R3615 VSS.n1383 VSS.t9 17.1921
R3616 VSS.n2627 VSS.n17 16.9417
R3617 VSS.n1058 VSS.n1057 16.9417
R3618 VSS.n1356 VSS.n718 16.6711
R3619 VSS.n1363 VSS.n713 16.6711
R3620 VSS.n1365 VSS.n1364 16.6711
R3621 VSS.n1419 VSS.n1418 16.6711
R3622 VSS.n903 VSS.n702 16.6711
R3623 VSS.n1412 VSS.n708 16.6711
R3624 VSS.n1411 VSS.n1376 16.6711
R3625 VSS.n1379 VSS.n1378 16.6711
R3626 VSS.n1644 VSS.n507 16.6711
R3627 VSS.t30 VSS.n718 16.1502
R3628 VSS.n671 VSS.n665 15.8123
R3629 VSS.n1461 VSS.n1435 15.8123
R3630 VSS.n811 VSS.n810 15.8123
R3631 VSS.n870 VSS.n842 15.8123
R3632 VSS.n1628 VSS.n571 15.6292
R3633 VSS.n1622 VSS.n1621 15.6292
R3634 VSS.n585 VSS.n578 15.6292
R3635 VSS.n1615 VSS.n586 15.6292
R3636 VSS.n993 VSS.n593 15.6292
R3637 VSS.n1608 VSS.n1607 15.6292
R3638 VSS.n1001 VSS.n595 15.6292
R3639 VSS.n1600 VSS.n602 15.6292
R3640 VSS.n1550 VSS.n1549 15.6292
R3641 VSS.n2100 VSS.t34 15.1082
R3642 VSS.t38 VSS.n2029 15.1082
R3643 VSS.n1593 VSS.n608 15.1082
R3644 VSS.n478 VSS.n477 14.5711
R3645 VSS.n463 VSS.n457 14.5711
R3646 VSS.n437 VSS.n436 14.5711
R3647 VSS.n417 VSS.n409 14.5711
R3648 VSS.n1686 VSS.n1675 14.5711
R3649 VSS.n1690 VSS.n1689 14.5711
R3650 VSS.n1673 VSS.n1672 14.5711
R3651 VSS.n1750 VSS.n1749 14.5711
R3652 VSS.n1746 VSS.n1735 14.5711
R3653 VSS.n1728 VSS.n1727 14.5711
R3654 VSS.n670 VSS.n667 14.3064
R3655 VSS.n1465 VSS.n1464 14.3064
R3656 VSS.n807 VSS.n805 14.3064
R3657 VSS.n872 VSS.n871 14.3064
R3658 VSS.n1369 VSS.n1368 14.3064
R3659 VSS.t14 VSS.n2068 14.0663
R3660 VSS.n2061 VSS.t26 14.0663
R3661 VSS.n778 VSS.n770 13.9299
R3662 VSS.n2361 VSS.n2360 13.9299
R3663 VSS.n1350 VSS.n1349 13.9299
R3664 VSS.n2550 VSS.n2549 13.9299
R3665 VSS.n28 VSS.n15 13.5534
R3666 VSS.n1053 VSS.n997 13.5534
R3667 VSS.t8 VSS.n569 13.5454
R3668 VSS.n2628 VSS.n2627 13.177
R3669 VSS.n1057 VSS.n1056 13.177
R3670 VSS.n2315 VSS.n139 13.177
R3671 VSS.n253 VSS.t5 13.0244
R3672 VSS.n2022 VSS.t0 13.0244
R3673 VSS.n1494 VSS.t60 13.0244
R3674 VSS.n1494 VSS.n1493 12.5035
R3675 VSS.n644 VSS.n643 12.5035
R3676 VSS.n643 VSS.t13 12.5035
R3677 VSS.n2557 VSS.n2556 12.5035
R3678 VSS.n59 VSS.n57 12.5035
R3679 VSS.n2563 VSS.n52 12.5035
R3680 VSS.n2547 VSS.n2546 12.5035
R3681 VSS.n2628 VSS.n18 12.424
R3682 VSS.n1056 VSS.n995 12.424
R3683 VSS.n146 VSS.n139 12.424
R3684 VSS.n26 VSS.n15 12.0476
R3685 VSS.n1053 VSS.n1052 12.0476
R3686 VSS.n1637 VSS.n513 11.9825
R3687 VSS.n1614 VSS.t22 11.9825
R3688 VSS.n778 VSS.n777 11.6711
R3689 VSS.n2360 VSS.n117 11.6711
R3690 VSS.n1354 VSS.n1350 11.6711
R3691 VSS.n2550 VSS.n62 11.6711
R3692 VSS.n671 VSS.n670 11.2946
R3693 VSS.n1464 VSS.n1435 11.2946
R3694 VSS.n810 VSS.n805 11.2946
R3695 VSS.n871 VSS.n870 11.2946
R3696 VSS.n1369 VSS.n710 11.2946
R3697 VSS.n1472 VSS.n1471 11.0636
R3698 VSS.n1470 VSS.n692 11.0636
R3699 VSS.n1469 VSS.n693 11.0636
R3700 VSS.n1468 VSS.n1467 11.0636
R3701 VSS.n1473 VSS.n691 11.0636
R3702 VSS.n1475 VSS.n1474 11.0636
R3703 VSS.n1477 VSS.n1476 11.0636
R3704 VSS.n1478 VSS.n655 11.0636
R3705 VSS.n1480 VSS.n1479 11.0636
R3706 VSS.n879 VSS.n835 11.0636
R3707 VSS.n834 VSS.n792 11.0636
R3708 VSS.n833 VSS.n793 11.0636
R3709 VSS.n832 VSS.n794 11.0636
R3710 VSS.n831 VSS.n830 11.0636
R3711 VSS.n878 VSS.n836 11.0636
R3712 VSS.n877 VSS.n837 11.0636
R3713 VSS.n876 VSS.n838 11.0636
R3714 VSS.n875 VSS.n874 11.0636
R3715 VSS.t8 VSS.n563 10.9406
R3716 VSS.n1630 VSS.n569 10.9406
R3717 VSS.n1357 VSS.t57 10.4196
R3718 VSS.t7 VSS.n1376 10.4196
R3719 VSS.n1622 VSS.t23 10.4196
R3720 VSS.n2557 VSS.t13 10.4196
R3721 VSS.n45 VSS.t59 10.4196
R3722 VSS.t33 VSS.n886 10.2467
R3723 VSS.n1020 VSS.t22 10.2467
R3724 VSS.t43 VSS.n708 9.89868
R3725 VSS.n645 VSS.t60 9.89868
R3726 VSS.n674 VSS.n665 9.78874
R3727 VSS.n1461 VSS.n1460 9.78874
R3728 VSS.n811 VSS.n803 9.78874
R3729 VSS.n867 VSS.n842 9.78874
R3730 VSS.n689 VSS.n657 9.58499
R3731 VSS.n1445 VSS.n1444 9.58499
R3732 VSS.n827 VSS.n795 9.58499
R3733 VSS.n851 VSS.n850 9.58499
R3734 VSS.n2310 VSS.n137 9.52595
R3735 VSS.n2551 VSS.n2550 9.49023
R3736 VSS.n1488 VSS.n650 9.49023
R3737 VSS.n1391 VSS.n598 9.49023
R3738 VSS.n1400 VSS.n1396 9.49023
R3739 VSS.n1026 VSS.n1015 9.49023
R3740 VSS.n928 VSS.n783 9.49023
R3741 VSS.n1031 VSS.n1013 9.49023
R3742 VSS.n2360 VSS.n2359 9.49023
R3743 VSS.n909 VSS.n908 9.49023
R3744 VSS.n779 VSS.n778 9.49023
R3745 VSS.n1972 VSS.n1971 9.49023
R3746 VSS.n1797 VSS.n399 9.49023
R3747 VSS.n1352 VSS.n1350 9.49023
R3748 VSS.n1408 VSS.n1407 9.49023
R3749 VSS.n2603 VSS.n14 9.41955
R3750 VSS.n2629 VSS.n17 9.41955
R3751 VSS.n1065 VSS.n1064 9.41955
R3752 VSS.n1370 VSS.n1369 9.41955
R3753 VSS.n998 VSS.n996 9.35854
R3754 VSS.n657 VSS.n656 9.3005
R3755 VSS.n686 VSS.n685 9.3005
R3756 VSS.n684 VSS.n683 9.3005
R3757 VSS.n661 VSS.n660 9.3005
R3758 VSS.n678 VSS.n677 9.3005
R3759 VSS.n676 VSS.n675 9.3005
R3760 VSS.n665 VSS.n664 9.3005
R3761 VSS.n670 VSS.n669 9.3005
R3762 VSS.n1446 VSS.n1445 9.3005
R3763 VSS.n1448 VSS.n1447 9.3005
R3764 VSS.n1441 VSS.n1440 9.3005
R3765 VSS.n1454 VSS.n1453 9.3005
R3766 VSS.n1456 VSS.n1455 9.3005
R3767 VSS.n1437 VSS.n1436 9.3005
R3768 VSS.n1462 VSS.n1461 9.3005
R3769 VSS.n1464 VSS.n1463 9.3005
R3770 VSS.n828 VSS.n827 9.3005
R3771 VSS.n797 VSS.n796 9.3005
R3772 VSS.n822 VSS.n821 9.3005
R3773 VSS.n820 VSS.n819 9.3005
R3774 VSS.n801 VSS.n800 9.3005
R3775 VSS.n814 VSS.n813 9.3005
R3776 VSS.n812 VSS.n811 9.3005
R3777 VSS.n805 VSS.n804 9.3005
R3778 VSS.n850 VSS.n849 9.3005
R3779 VSS.n855 VSS.n854 9.3005
R3780 VSS.n857 VSS.n856 9.3005
R3781 VSS.n846 VSS.n845 9.3005
R3782 VSS.n863 VSS.n862 9.3005
R3783 VSS.n866 VSS.n865 9.3005
R3784 VSS.n864 VSS.n842 9.3005
R3785 VSS.n871 VSS.n841 9.3005
R3786 VSS.n2608 VSS.n14 9.3005
R3787 VSS.n2630 VSS.n16 9.3005
R3788 VSS.n2630 VSS.n15 9.3005
R3789 VSS.n2629 VSS.n2628 9.3005
R3790 VSS.n460 VSS.n459 9.3005
R3791 VSS.n462 VSS.n461 9.3005
R3792 VSS.n472 VSS.n471 9.3005
R3793 VSS.n474 VSS.n473 9.3005
R3794 VSS.n451 VSS.n450 9.3005
R3795 VSS.n425 VSS.n415 9.3005
R3796 VSS.n418 VSS.n416 9.3005
R3797 VSS.n420 VSS.n419 9.3005
R3798 VSS.n433 VSS.n432 9.3005
R3799 VSS.n411 VSS.n410 9.3005
R3800 VSS.n1677 VSS.n1676 9.3005
R3801 VSS.n1655 VSS.n1654 9.3005
R3802 VSS.n1669 VSS.n1668 9.3005
R3803 VSS.n1667 VSS.n1666 9.3005
R3804 VSS.n1661 VSS.n1660 9.3005
R3805 VSS.n1683 VSS.n1682 9.3005
R3806 VSS.n1685 VSS.n1684 9.3005
R3807 VSS.n1743 VSS.n1742 9.3005
R3808 VSS.n1745 VSS.n1744 9.3005
R3809 VSS.n1724 VSS.n1723 9.3005
R3810 VSS.n1722 VSS.n1721 9.3005
R3811 VSS.n1716 VSS.n1715 9.3005
R3812 VSS.n1738 VSS.n1737 9.3005
R3813 VSS.n1730 VSS.n1729 9.3005
R3814 VSS.n361 VSS.n359 9.3005
R3815 VSS.n1960 VSS.n1959 9.3005
R3816 VSS.n353 VSS.n352 9.3005
R3817 VSS.n1971 VSS.n1970 9.3005
R3818 VSS.n358 VSS.n355 9.3005
R3819 VSS.n1958 VSS.n1957 9.3005
R3820 VSS.n1949 VSS.n363 9.3005
R3821 VSS.n1787 VSS.n1786 9.3005
R3822 VSS.n1796 VSS.n1795 9.3005
R3823 VSS.n1785 VSS.n1784 9.3005
R3824 VSS.n402 VSS.n401 9.3005
R3825 VSS.n1798 VSS.n1797 9.3005
R3826 VSS.n408 VSS.n404 9.3005
R3827 VSS.n1779 VSS.n1753 9.3005
R3828 VSS.n1056 VSS.n1055 9.3005
R3829 VSS.n1054 VSS.n1053 9.3005
R3830 VSS.n1058 VSS.n991 9.3005
R3831 VSS.n1064 VSS.n1063 9.3005
R3832 VSS.n1371 VSS.n1370 9.3005
R3833 VSS.n1373 VSS.n502 9.3005
R3834 VSS.n1648 VSS.n1647 9.3005
R3835 VSS.n139 VSS.n137 9.3005
R3836 VSS.n2317 VSS.n2316 9.3005
R3837 VSS.n779 VSS.n774 9.3005
R3838 VSS.n1084 VSS.n1083 9.3005
R3839 VSS.n908 VSS.n907 9.3005
R3840 VSS.n930 VSS.n783 9.3005
R3841 VSS.n1076 VSS.n1075 9.3005
R3842 VSS.n1026 VSS.n1025 9.3005
R3843 VSS.n1032 VSS.n1031 9.3005
R3844 VSS.n2350 VSS.n2349 9.3005
R3845 VSS.n2359 VSS.n2358 9.3005
R3846 VSS.n1400 VSS.n1399 9.3005
R3847 VSS.n2552 VSS.n2551 9.3005
R3848 VSS.n1482 VSS.n61 9.3005
R3849 VSS.n1489 VSS.n1488 9.3005
R3850 VSS.n1391 VSS.n1390 9.3005
R3851 VSS.n1618 VSS.n582 9.3005
R3852 VSS.n1353 VSS.n1352 9.3005
R3853 VSS.n1423 VSS.n1422 9.3005
R3854 VSS.n1407 VSS.n1406 9.3005
R3855 VSS.t43 VSS.n903 8.85676
R3856 VSS.n2579 VSS.n17 8.65932
R3857 VSS.n1059 VSS.n1058 8.65932
R3858 VSS.n1379 VSS.t7 8.33581
R3859 VSS.n1069 VSS.n1068 8.33581
R3860 VSS.n675 VSS.n663 8.28285
R3861 VSS.n1457 VSS.n1437 8.28285
R3862 VSS.n815 VSS.n814 8.28285
R3863 VSS.n866 VSS.n844 8.28285
R3864 VSS.n1970 VSS.n351 8.28285
R3865 VSS.n1799 VSS.n1798 8.28285
R3866 VSS.n1063 VSS.n990 8.28285
R3867 VSS.n1670 VSS.n1665 8.2073
R3868 VSS.n1725 VSS.n1720 8.2073
R3869 VSS.n2092 VSS.t16 7.81485
R3870 VSS.t20 VSS.n2037 7.81485
R3871 VSS.n1541 VSS.n624 7.81485
R3872 VSS.n2604 VSS.n16 7.52991
R3873 VSS.n1000 VSS.n998 7.52991
R3874 VSS.t30 VSS.n1088 7.3192
R3875 VSS.n2355 VSS.t2 7.3192
R3876 VSS.n1070 VSS.n1069 7.29389
R3877 VSS.n199 VSS.n198 7.24494
R3878 VSS.n2609 VSS.n2608 7.15344
R3879 VSS.n931 VSS.n928 7.15344
R3880 VSS.n1024 VSS.n1015 7.15344
R3881 VSS.n1398 VSS.n1396 7.15344
R3882 VSS.n1389 VSS.n598 7.15344
R3883 VSS.n679 VSS.n678 6.77697
R3884 VSS.n1456 VSS.n1439 6.77697
R3885 VSS.n818 VSS.n801 6.77697
R3886 VSS.n862 VSS.n861 6.77697
R3887 VSS.n1372 VSS.n1371 6.77697
R3888 VSS.t55 VSS.n2076 6.77294
R3889 VSS.n2053 VSS.t3 6.77294
R3890 VSS.n458 VSS.n455 6.41949
R3891 VSS.n431 VSS.n412 6.41949
R3892 VSS.n1681 VSS.n1658 6.41949
R3893 VSS.n1678 VSS.n1656 6.41949
R3894 VSS.n1739 VSS.n1731 6.41949
R3895 VSS.n1741 VSS.n1733 6.41949
R3896 VSS.n1277 VSS.t57 6.25198
R3897 VSS.n464 VSS.t135 5.8005
R3898 VSS.t92 VSS.n464 5.8005
R3899 VSS.n465 VSS.t92 5.8005
R3900 VSS.n465 VSS.t115 5.8005
R3901 VSS.n447 VSS.t40 5.8005
R3902 VSS.n447 VSS.t62 5.8005
R3903 VSS.n445 VSS.t47 5.8005
R3904 VSS.n445 VSS.t29 5.8005
R3905 VSS.n443 VSS.t15 5.8005
R3906 VSS.n443 VSS.t46 5.8005
R3907 VSS.n441 VSS.t54 5.8005
R3908 VSS.n441 VSS.t61 5.8005
R3909 VSS.n439 VSS.t35 5.8005
R3910 VSS.n439 VSS.t63 5.8005
R3911 VSS.n435 VSS.t124 5.8005
R3912 VSS.n435 VSS.t41 5.8005
R3913 VSS.n428 VSS.t126 5.8005
R3914 VSS.n428 VSS.t124 5.8005
R3915 VSS.t128 VSS.n1687 5.8005
R3916 VSS.n1687 VSS.t85 5.8005
R3917 VSS.n1688 VSS.t137 5.8005
R3918 VSS.n1688 VSS.t128 5.8005
R3919 VSS.n1671 VSS.t136 5.8005
R3920 VSS.n1671 VSS.t78 5.8005
R3921 VSS.n1748 VSS.t96 5.8005
R3922 VSS.n1748 VSS.t94 5.8005
R3923 VSS.t94 VSS.n1747 5.8005
R3924 VSS.n1747 VSS.t44 5.8005
R3925 VSS.n1726 VSS.t89 5.8005
R3926 VSS.n1726 VSS.t37 5.8005
R3927 VSS.n1692 VSS.t42 5.8005
R3928 VSS.n1692 VSS.t1 5.8005
R3929 VSS.n1696 VSS.t25 5.8005
R3930 VSS.n1696 VSS.t133 5.8005
R3931 VSS.n1700 VSS.t31 5.8005
R3932 VSS.n1700 VSS.t4 5.8005
R3933 VSS.n1704 VSS.t134 5.8005
R3934 VSS.n1704 VSS.t58 5.8005
R3935 VSS.n1708 VSS.t32 5.8005
R3936 VSS.n1708 VSS.t138 5.8005
R3937 VSS.n1712 VSS.t6 5.8005
R3938 VSS.n1712 VSS.t45 5.8005
R3939 VSS.n1694 VSS.t21 5.8005
R3940 VSS.n1694 VSS.t39 5.8005
R3941 VSS.n1698 VSS.t28 5.8005
R3942 VSS.n1698 VSS.t51 5.8005
R3943 VSS.n1702 VSS.t48 5.8005
R3944 VSS.n1702 VSS.t27 5.8005
R3945 VSS.n1706 VSS.t64 5.8005
R3946 VSS.n1706 VSS.t56 5.8005
R3947 VSS.n1710 VSS.t50 5.8005
R3948 VSS.n1710 VSS.t17 5.8005
R3949 VSS.n246 VSS.t36 5.73102
R3950 VSS.n2014 VSS.t91 5.73102
R3951 VSS.t33 VSS.t23 5.73102
R3952 VSS.t11 VSS.t52 5.73102
R3953 VSS.n1960 VSS.n357 5.64756
R3954 VSS.n1787 VSS.n403 5.64756
R3955 VSS.n472 VSS.n468 5.37662
R3956 VSS.n427 VSS.n415 5.37662
R3957 VSS.n682 VSS.n661 5.27109
R3958 VSS.n1453 VSS.n1452 5.27109
R3959 VSS.n819 VSS.n799 5.27109
R3960 VSS.n858 VSS.n846 5.27109
R3961 VSS.n1086 VSS.n774 5.27109
R3962 VSS.n2358 VSS.n2357 5.27109
R3963 VSS.n1353 VSS.n1351 5.27109
R3964 VSS.n2553 VSS.n2552 5.27109
R3965 VSS.n1601 VSS.t52 5.21007
R3966 VSS.n2547 VSS.t19 5.21007
R3967 VSS.n2117 VSS.n239 4.68911
R3968 VSS.n1049 VSS.t11 4.68911
R3969 VSS.n1964 VSS.n355 4.51815
R3970 VSS.n1950 VSS.n361 4.51815
R3971 VSS.n1791 VSS.n402 4.51815
R3972 VSS.n1780 VSS.n408 4.51815
R3973 VSS.n1084 VSS.n775 4.51815
R3974 VSS.n2351 VSS.n2350 4.51815
R3975 VSS.n1422 VSS.n1421 4.51815
R3976 VSS.n1490 VSS.n61 4.51815
R3977 VSS.n2346 VSS.n118 4.5005
R3978 VSS.n1030 VSS.n1029 4.5005
R3979 VSS.n128 VSS.n127 4.5005
R3980 VSS.n2348 VSS.n2347 4.5005
R3981 VSS.n1079 VSS.n1078 4.5005
R3982 VSS.n1077 VSS.n782 4.5005
R3983 VSS.n1014 VSS.n881 4.5005
R3984 VSS.n1028 VSS.n1027 4.5005
R3985 VSS.n1080 VSS.n781 4.5005
R3986 VSS.n1082 VSS.n1081 4.5005
R3987 VSS.n1405 VSS.n1404 4.5005
R3988 VSS.n1388 VSS.n696 4.5005
R3989 VSS.n1392 VSS.n652 4.5005
R3990 VSS.n1403 VSS.n1402 4.5005
R3991 VSS.n1401 VSS.n1395 4.5005
R3992 VSS.n1394 VSS.n1393 4.5005
R3993 VSS.n653 VSS.n63 4.5005
R3994 VSS.n1484 VSS.n1483 4.5005
R3995 VSS.n1485 VSS.n651 4.5005
R3996 VSS.n1487 VSS.n1486 4.5005
R3997 VSS.n1651 VSS.n479 4.26732
R3998 VSS.n1345 VSS.n1344 4.16815
R3999 VSS.n438 VSS.n409 3.81995
R4000 VSS.n683 VSS.n659 3.76521
R4001 VSS.n1449 VSS.n1441 3.76521
R4002 VSS.n823 VSS.n822 3.76521
R4003 VSS.n857 VSS.n848 3.76521
R4004 VSS.n475 VSS.n451 3.76521
R4005 VSS.n462 VSS.n456 3.76521
R4006 VSS.n434 VSS.n411 3.76521
R4007 VSS.n421 VSS.n420 3.76521
R4008 VSS.n1685 VSS.n1659 3.76521
R4009 VSS.n1657 VSS.n1655 3.76521
R4010 VSS.n1662 VSS.n1661 3.76521
R4011 VSS.n1732 VSS.n1730 3.76521
R4012 VSS.n1745 VSS.n1734 3.76521
R4013 VSS.n1717 VSS.n1716 3.76521
R4014 VSS.n1066 VSS.n1065 3.76521
R4015 VSS.n1374 VSS.n1373 3.76521
R4016 VSS.n907 VSS.n898 3.76521
R4017 VSS.n1033 VSS.n1032 3.76521
R4018 VSS.n1406 VSS.n1381 3.76521
R4019 VSS.n1489 VSS.n647 3.76521
R4020 VSS.n2318 VSS.n2317 3.68738
R4021 VSS.t33 VSS.n1070 3.6472
R4022 VSS.n992 VSS.t22 3.6472
R4023 VSS.n1651 VSS.n1650 3.44797
R4024 VSS.n2343 VSS.n129 3.4105
R4025 VSS.n2638 VSS.n2637 3.4105
R4026 VSS.n2643 VSS.n8 3.4105
R4027 VSS.n497 VSS.n496 3.4105
R4028 VSS.n489 VSS.n485 3.4105
R4029 VSS.n132 VSS.n131 3.4105
R4030 VSS.n2320 VSS.n136 3.4105
R4031 VSS.n2654 VSS.n3 3.4105
R4032 VSS.n2650 VSS.n2649 3.4105
R4033 VSS.n2654 VSS.n1 3.4105
R4034 VSS.n2338 VSS.n2334 3.4105
R4035 VSS.n2343 VSS.n2342 3.4105
R4036 VSS.n485 VSS.n484 3.4105
R4037 VSS.n2639 VSS.n2638 3.4105
R4038 VSS.n2643 VSS.n6 3.4105
R4039 VSS.n131 VSS.n130 3.4105
R4040 VSS.n669 VSS.n668 3.09986
R4041 VSS.n1463 VSS.n1433 3.09986
R4042 VSS.n806 VSS.n804 3.09986
R4043 VSS.n873 VSS.n841 3.09986
R4044 VSS.n1691 VSS.n1690 2.89851
R4045 VSS.n1735 VSS.n1714 2.89851
R4046 VSS.n501 VSS.n500 2.72553
R4047 VSS.n457 VSS.n449 2.67025
R4048 VSS.n479 VSS.n478 2.67025
R4049 VSS.n438 VSS.n437 2.67025
R4050 VSS.n2612 VSS.n2603 2.63579
R4051 VSS.n910 VSS.n909 2.63579
R4052 VSS.n1034 VSS.n1013 2.63579
R4053 VSS.n1409 VSS.n1408 2.63579
R4054 VSS.n650 VSS.n649 2.63579
R4055 VSS.t30 VSS.n713 2.60528
R4056 VSS.n59 VSS.t2 2.60528
R4057 VSS.n1473 VSS.t108 2.48621
R4058 VSS.t106 VSS.n1473 2.48621
R4059 VSS.n1472 VSS.t132 2.48621
R4060 VSS.t108 VSS.n1472 2.48621
R4061 VSS.t66 VSS.n692 2.48621
R4062 VSS.n692 VSS.t132 2.48621
R4063 VSS.t70 VSS.n693 2.48621
R4064 VSS.n693 VSS.t66 2.48621
R4065 VSS.n1467 VSS.t75 2.48621
R4066 VSS.n1467 VSS.t70 2.48621
R4067 VSS.n1474 VSS.t106 2.48621
R4068 VSS.n1474 VSS.t102 2.48621
R4069 VSS.n1477 VSS.t102 2.48621
R4070 VSS.t100 VSS.n1477 2.48621
R4071 VSS.n1478 VSS.t100 2.48621
R4072 VSS.t120 VSS.n1478 2.48621
R4073 VSS.n1479 VSS.t120 2.48621
R4074 VSS.n1479 VSS.t72 2.48621
R4075 VSS.t118 VSS.n835 2.48621
R4076 VSS.n835 VSS.t130 2.48621
R4077 VSS.t130 VSS.n834 2.48621
R4078 VSS.n834 VSS.t81 2.48621
R4079 VSS.t81 VSS.n833 2.48621
R4080 VSS.n833 VSS.t98 2.48621
R4081 VSS.t98 VSS.n832 2.48621
R4082 VSS.n832 VSS.t113 2.48621
R4083 VSS.t113 VSS.n831 2.48621
R4084 VSS.n831 VSS.t110 2.48621
R4085 VSS.t122 VSS.n836 2.48621
R4086 VSS.n836 VSS.t118 2.48621
R4087 VSS.t104 VSS.n837 2.48621
R4088 VSS.n837 VSS.t122 2.48621
R4089 VSS.t83 VSS.n838 2.48621
R4090 VSS.n838 VSS.t104 2.48621
R4091 VSS.n874 VSS.t68 2.48621
R4092 VSS.n874 VSS.t83 2.48621
R4093 VSS.n1081 VSS.n780 2.30235
R4094 VSS.n1388 VSS.n695 2.30235
R4095 VSS.n2636 VSS.n2635 2.27039
R4096 VSS.n2321 VSS.n2318 2.27036
R4097 VSS.n500 VSS.n480 2.27013
R4098 VSS.n687 VSS.n686 2.25932
R4099 VSS.n1448 VSS.n1443 2.25932
R4100 VSS.n826 VSS.n797 2.25932
R4101 VSS.n854 VSS.n853 2.25932
R4102 VSS.n474 VSS.n453 2.25932
R4103 VSS.n424 VSS.n416 2.25932
R4104 VSS.n1666 VSS.n1663 2.25932
R4105 VSS.n1721 VSS.n1718 2.25932
R4106 VSS.n1674 VSS.n1653 2.25177
R4107 VSS.n1752 VSS.n1751 2.25177
R4108 VSS.n2633 VSS.n2632 2.2505
R4109 VSS.n490 VSS.n481 2.2505
R4110 VSS.n2328 VSS.n2327 2.2505
R4111 VSS.t12 VSS.n992 2.08433
R4112 VSS.n1593 VSS.t10 2.08433
R4113 VSS.n2346 VSS.n2345 2.0166
R4114 VSS.n653 VSS.n2 2.0166
R4115 VSS.n1029 VSS.n1028 2.00152
R4116 VSS.n1080 VSS.n1079 2.00152
R4117 VSS.n1404 VSS.n1403 2.00152
R4118 VSS.n1486 VSS.n652 2.00152
R4119 VSS.n1648 VSS.n503 1.94348
R4120 VSS.n1973 VSS.n1972 1.88285
R4121 VSS.n1965 VSS.n353 1.88285
R4122 VSS.n1802 VSS.n399 1.88285
R4123 VSS.n1795 VSS.n1794 1.88285
R4124 VSS.n1753 VSS.n1752 1.82131
R4125 VSS.n1650 VSS.n501 1.74238
R4126 VSS.n2644 VSS.n7 1.71461
R4127 VSS.n488 VSS.n487 1.71461
R4128 VSS.n2330 VSS.n2329 1.71461
R4129 VSS.n2337 VSS.n0 1.70929
R4130 VSS.n2648 VSS.n2646 1.70929
R4131 VSS.n495 VSS.n480 1.70926
R4132 VSS.n2322 VSS.n2321 1.70926
R4133 VSS.n2345 VSS.n2344 1.7055
R4134 VSS.n2335 VSS.n2333 1.7055
R4135 VSS.n2339 VSS.n2336 1.7055
R4136 VSS.n2642 VSS.n9 1.7055
R4137 VSS.n2631 VSS.n10 1.7055
R4138 VSS.n2636 VSS.n12 1.7055
R4139 VSS.n492 VSS.n491 1.7055
R4140 VSS.n483 VSS.n482 1.7055
R4141 VSS.n135 VSS.n134 1.7055
R4142 VSS.n2326 VSS.n2325 1.7055
R4143 VSS.n2655 VSS.n2 1.7055
R4144 VSS.n2653 VSS.n4 1.7055
R4145 VSS.n2647 VSS.n5 1.7055
R4146 VSS.n2653 VSS.n2652 1.7055
R4147 VSS.n2656 VSS.n2655 1.7055
R4148 VSS.n2651 VSS.n5 1.7055
R4149 VSS.n2341 VSS.n2333 1.7055
R4150 VSS.n2344 VSS.n2332 1.7055
R4151 VSS.n2340 VSS.n2339 1.7055
R4152 VSS.n493 VSS.n492 1.7055
R4153 VSS.n487 VSS.n486 1.7055
R4154 VSS.n494 VSS.n483 1.7055
R4155 VSS.n2642 VSS.n2641 1.7055
R4156 VSS.n2645 VSS.n2644 1.7055
R4157 VSS.n2640 VSS.n10 1.7055
R4158 VSS.n12 VSS.n11 1.7055
R4159 VSS.n2323 VSS.n135 1.7055
R4160 VSS.n2331 VSS.n2330 1.7055
R4161 VSS.n2325 VSS.n2324 1.7055
R4162 VSS.n1838 VSS.t88 1.56337
R4163 VSS.n2006 VSS.t77 1.56337
R4164 VSS.n1644 VSS.t9 1.56337
R4165 VSS.n1652 VSS.n363 1.20384
R4166 VSS.n2633 VSS.n7 1.20242
R4167 VSS.n488 VSS.n481 1.20242
R4168 VSS.n2329 VSS.n2328 1.20242
R4169 VSS.n2337 VSS.n2336 1.17304
R4170 VSS.n2648 VSS.n2647 1.17304
R4171 VSS.n440 VSS.n438 1.1502
R4172 VSS.n442 VSS.n440 1.1502
R4173 VSS.n444 VSS.n442 1.1502
R4174 VSS.n446 VSS.n444 1.1502
R4175 VSS.n448 VSS.n446 1.1502
R4176 VSS.n449 VSS.n448 1.1502
R4177 VSS.n479 VSS.n449 1.1502
R4178 VSS.n2323 VSS.n2322 1.14372
R4179 VSS.n495 VSS.n494 1.14372
R4180 VSS.n2634 VSS.n13 1.1255
R4181 VSS.n499 VSS.n498 1.1255
R4182 VSS.n2319 VSS.n133 1.1255
R4183 VSS.n1419 VSS.t18 1.04241
R4184 VSS.n1652 VSS.n1651 0.950967
R4185 VSS.n1471 VSS.n691 0.779912
R4186 VSS.n1471 VSS.n1470 0.779912
R4187 VSS.n1470 VSS.n1469 0.779912
R4188 VSS.n1468 VSS.n694 0.779912
R4189 VSS.n1469 VSS.n1468 0.779912
R4190 VSS.n1475 VSS.n691 0.779912
R4191 VSS.n1476 VSS.n1475 0.779912
R4192 VSS.n1476 VSS.n655 0.779912
R4193 VSS.n1480 VSS.n655 0.779912
R4194 VSS.n1480 VSS.n690 0.779912
R4195 VSS.n879 VSS.n792 0.779912
R4196 VSS.n793 VSS.n792 0.779912
R4197 VSS.n794 VSS.n793 0.779912
R4198 VSS.n830 VSS.n794 0.779912
R4199 VSS.n830 VSS.n829 0.779912
R4200 VSS.n879 VSS.n878 0.779912
R4201 VSS.n878 VSS.n877 0.779912
R4202 VSS.n877 VSS.n876 0.779912
R4203 VSS.n875 VSS.n839 0.779912
R4204 VSS.n876 VSS.n875 0.779912
R4205 VSS VSS.n0 0.765176
R4206 VSS.n471 VSS.n470 0.753441
R4207 VSS.n426 VSS.n425 0.753441
R4208 VSS.n1957 VSS.n360 0.753441
R4209 VSS.n1784 VSS.n407 0.753441
R4210 VSS.n1647 VSS.n504 0.753441
R4211 VSS.n930 VSS.n929 0.753441
R4212 VSS.n1025 VSS.n1016 0.753441
R4213 VSS.n1399 VSS.n581 0.753441
R4214 VSS.n1390 VSS.n583 0.753441
R4215 VSS.n1426 VSS.n1425 0.701719
R4216 VSS.n1425 VSS.n1424 0.701719
R4217 VSS.n1424 VSS.n654 0.701719
R4218 VSS.n1431 VSS.n1430 0.701719
R4219 VSS.n1430 VSS.n1429 0.701719
R4220 VSS.n1429 VSS.n1428 0.701719
R4221 VSS.n787 VSS.n786 0.701719
R4222 VSS.n786 VSS.n785 0.701719
R4223 VSS.n785 VSS.n784 0.701719
R4224 VSS.n789 VSS.n788 0.701719
R4225 VSS.n790 VSS.n789 0.701719
R4226 VSS.n791 VSS.n790 0.701719
R4227 VSS.n1675 VSS.n1674 0.647239
R4228 VSS.n1751 VSS.n1750 0.647239
R4229 VSS.n1653 VSS.n1652 0.617976
R4230 VSS.n1752 VSS.n1714 0.574311
R4231 VSS.n1714 VSS.n1713 0.574311
R4232 VSS.n1713 VSS.n1711 0.574311
R4233 VSS.n1711 VSS.n1709 0.574311
R4234 VSS.n1709 VSS.n1707 0.574311
R4235 VSS.n1707 VSS.n1705 0.574311
R4236 VSS.n1705 VSS.n1703 0.574311
R4237 VSS.n1703 VSS.n1701 0.574311
R4238 VSS.n1701 VSS.n1699 0.574311
R4239 VSS.n1699 VSS.n1697 0.574311
R4240 VSS.n1697 VSS.n1695 0.574311
R4241 VSS.n1695 VSS.n1693 0.574311
R4242 VSS.n1693 VSS.n1691 0.574311
R4243 VSS.n1691 VSS.n1653 0.574311
R4244 VSS.n2084 VSS.t53 0.521457
R4245 VSS.t24 VSS.n2045 0.521457
R4246 VSS.n1674 VSS.n1673 0.418978
R4247 VSS.n1751 VSS.n1728 0.418978
R4248 VSS.n458 VSS.n454 0.320353
R4249 VSS.n466 VSS.n454 0.320353
R4250 VSS.n467 VSS.n466 0.320353
R4251 VSS.n472 VSS.n467 0.320353
R4252 VSS.n415 VSS.n413 0.320353
R4253 VSS.n429 VSS.n413 0.320353
R4254 VSS.n430 VSS.n429 0.320353
R4255 VSS.n431 VSS.n430 0.320353
R4256 VSS.n1679 VSS.n1678 0.320353
R4257 VSS.n1681 VSS.n1679 0.320353
R4258 VSS.n1681 VSS.n1680 0.320353
R4259 VSS.n1665 VSS.n1664 0.320353
R4260 VSS.n1741 VSS.n1740 0.320353
R4261 VSS.n1739 VSS.n1736 0.320353
R4262 VSS.n1740 VSS.n1739 0.320353
R4263 VSS.n1720 VSS.n1719 0.320353
R4264 VSS.n996 VSS.n501 0.303278
R4265 VSS.n1650 VSS.n1649 0.303278
R4266 VSS.n1468 VSS.n1432 0.272321
R4267 VSS.n1427 VSS.n691 0.272321
R4268 VSS.n1481 VSS.n1480 0.272321
R4269 VSS.n830 VSS.n126 0.272321
R4270 VSS.n880 VSS.n879 0.272321
R4271 VSS.n875 VSS.n776 0.272321
R4272 VSS.n1427 VSS.n1426 0.261436
R4273 VSS.n1481 VSS.n654 0.261436
R4274 VSS.n1432 VSS.n1431 0.261436
R4275 VSS.n1428 VSS.n1427 0.261436
R4276 VSS.n880 VSS.n787 0.261436
R4277 VSS.n784 VSS.n126 0.261436
R4278 VSS.n788 VSS.n776 0.261436
R4279 VSS.n880 VSS.n791 0.261436
R4280 VSS.n1971 VSS.n352 0.243804
R4281 VSS.n1959 VSS.n358 0.243804
R4282 VSS.n1797 VSS.n1796 0.243804
R4283 VSS.n1786 VSS.n401 0.243804
R4284 VSS.n2317 VSS.n137 0.21925
R4285 VSS.n1958 VSS.n359 0.204927
R4286 VSS.n1785 VSS.n404 0.204927
R4287 VSS.n1064 VSS.n991 0.204369
R4288 VSS.n1055 VSS.n1054 0.204369
R4289 VSS.n669 VSS.n664 0.196152
R4290 VSS.n676 VSS.n664 0.196152
R4291 VSS.n677 VSS.n676 0.196152
R4292 VSS.n677 VSS.n660 0.196152
R4293 VSS.n684 VSS.n660 0.196152
R4294 VSS.n685 VSS.n684 0.196152
R4295 VSS.n685 VSS.n656 0.196152
R4296 VSS.n690 VSS.n656 0.196152
R4297 VSS.n1463 VSS.n1462 0.196152
R4298 VSS.n1462 VSS.n1436 0.196152
R4299 VSS.n1455 VSS.n1436 0.196152
R4300 VSS.n1455 VSS.n1454 0.196152
R4301 VSS.n1454 VSS.n1440 0.196152
R4302 VSS.n1447 VSS.n1440 0.196152
R4303 VSS.n1447 VSS.n1446 0.196152
R4304 VSS.n1446 VSS.n694 0.196152
R4305 VSS.n829 VSS.n828 0.196152
R4306 VSS.n828 VSS.n796 0.196152
R4307 VSS.n821 VSS.n796 0.196152
R4308 VSS.n821 VSS.n820 0.196152
R4309 VSS.n820 VSS.n800 0.196152
R4310 VSS.n813 VSS.n800 0.196152
R4311 VSS.n813 VSS.n812 0.196152
R4312 VSS.n812 VSS.n804 0.196152
R4313 VSS.n849 VSS.n839 0.196152
R4314 VSS.n855 VSS.n849 0.196152
R4315 VSS.n856 VSS.n855 0.196152
R4316 VSS.n856 VSS.n845 0.196152
R4317 VSS.n863 VSS.n845 0.196152
R4318 VSS.n865 VSS.n863 0.196152
R4319 VSS.n865 VSS.n864 0.196152
R4320 VSS.n864 VSS.n841 0.196152
R4321 VSS.n461 VSS.n457 0.196152
R4322 VSS.n461 VSS.n460 0.196152
R4323 VSS.n460 VSS.n458 0.196152
R4324 VSS.n478 VSS.n450 0.196152
R4325 VSS.n473 VSS.n450 0.196152
R4326 VSS.n473 VSS.n472 0.196152
R4327 VSS.n419 VSS.n409 0.196152
R4328 VSS.n419 VSS.n418 0.196152
R4329 VSS.n418 VSS.n415 0.196152
R4330 VSS.n437 VSS.n410 0.196152
R4331 VSS.n432 VSS.n410 0.196152
R4332 VSS.n432 VSS.n431 0.196152
R4333 VSS.n1690 VSS.n1654 0.196152
R4334 VSS.n1677 VSS.n1654 0.196152
R4335 VSS.n1678 VSS.n1677 0.196152
R4336 VSS.n1668 VSS.n1665 0.196152
R4337 VSS.n1668 VSS.n1667 0.196152
R4338 VSS.n1667 VSS.n1660 0.196152
R4339 VSS.n1673 VSS.n1660 0.196152
R4340 VSS.n1684 VSS.n1675 0.196152
R4341 VSS.n1684 VSS.n1683 0.196152
R4342 VSS.n1683 VSS.n1681 0.196152
R4343 VSS.n1744 VSS.n1735 0.196152
R4344 VSS.n1744 VSS.n1743 0.196152
R4345 VSS.n1743 VSS.n1741 0.196152
R4346 VSS.n1723 VSS.n1720 0.196152
R4347 VSS.n1723 VSS.n1722 0.196152
R4348 VSS.n1722 VSS.n1715 0.196152
R4349 VSS.n1728 VSS.n1715 0.196152
R4350 VSS.n1750 VSS.n1729 0.196152
R4351 VSS.n1738 VSS.n1729 0.196152
R4352 VSS.n1739 VSS.n1738 0.196152
R4353 VSS.n358 VSS.n352 0.190232
R4354 VSS.n1959 VSS.n1958 0.190232
R4355 VSS.n1796 VSS.n401 0.190232
R4356 VSS.n1786 VSS.n1785 0.190232
R4357 VSS.n2646 VSS.n2645 0.181806
R4358 VSS.n2332 VSS.n2331 0.175397
R4359 VSS VSS.n2656 0.173973
R4360 VSS.n1483 VSS.n63 0.146333
R4361 VSS.n1487 VSS.n651 0.146333
R4362 VSS.n1393 VSS.n1392 0.146333
R4363 VSS.n1402 VSS.n1401 0.146333
R4364 VSS.n1027 VSS.n881 0.146333
R4365 VSS.n1078 VSS.n1077 0.146333
R4366 VSS.n1030 VSS.n127 0.146333
R4367 VSS.n2348 VSS.n118 0.146333
R4368 VSS.n1082 VSS.n781 0.146333
R4369 VSS.n1405 VSS.n696 0.146333
R4370 VSS.n780 VSS.n779 0.144812
R4371 VSS.n1352 VSS.n695 0.144812
R4372 VSS.n1083 VSS.n780 0.119763
R4373 VSS.n1423 VSS.n695 0.119763
R4374 VSS.n1055 VSS.n991 0.119548
R4375 VSS.n1432 VSS.n1423 0.114136
R4376 VSS.n1427 VSS.n582 0.114136
R4377 VSS.n1482 VSS.n1481 0.114136
R4378 VSS.n2349 VSS.n126 0.114136
R4379 VSS.n1076 VSS.n880 0.114136
R4380 VSS.n1083 VSS.n776 0.114136
R4381 VSS.n1370 VSS.n502 0.113595
R4382 VSS.n2635 VSS.n2630 0.113
R4383 VSS.n2630 VSS.n14 0.112107
R4384 VSS.n486 VSS.n11 0.110594
R4385 VSS.n363 VSS.n359 0.104667
R4386 VSS.n1753 VSS.n404 0.104667
R4387 VSS.n2630 VSS.n2629 0.0927619
R4388 VSS.n1029 VSS.n128 0.0788898
R4389 VSS.n2347 VSS.n2346 0.0788898
R4390 VSS.n1079 VSS.n782 0.0788898
R4391 VSS.n1028 VSS.n1014 0.0788898
R4392 VSS.n1081 VSS.n1080 0.0788898
R4393 VSS.n1404 VSS.n1388 0.0788898
R4394 VSS.n1403 VSS.n1395 0.0788898
R4395 VSS.n1394 VSS.n652 0.0788898
R4396 VSS.n1486 VSS.n1485 0.0788898
R4397 VSS.n1484 VSS.n653 0.0788898
R4398 VSS.n499 VSS.n481 0.0782244
R4399 VSS.n2551 VSS.n63 0.0719286
R4400 VSS.n1488 VSS.n1487 0.0719286
R4401 VSS.n1392 VSS.n1391 0.0719286
R4402 VSS.n1402 VSS.n1400 0.0719286
R4403 VSS.n1027 VSS.n1026 0.0719286
R4404 VSS.n1078 VSS.n783 0.0719286
R4405 VSS.n1031 VSS.n1030 0.0719286
R4406 VSS.n2359 VSS.n118 0.0719286
R4407 VSS.n908 VSS.n781 0.0719286
R4408 VSS.n1407 VSS.n1405 0.0719286
R4409 VSS.n2347 VSS.n128 0.0682966
R4410 VSS.n1014 VSS.n782 0.0682966
R4411 VSS.n1395 VSS.n1394 0.0682966
R4412 VSS.n1485 VSS.n1484 0.0682966
R4413 VSS.n2336 VSS.n2335 0.0675573
R4414 VSS.n2647 VSS.n4 0.0675573
R4415 VSS.n500 VSS.n499 0.0654412
R4416 VSS.n1054 VSS.n996 0.0615119
R4417 VSS.n1649 VSS.n502 0.0600238
R4418 VSS.n1649 VSS.n1648 0.0600238
R4419 VSS.n2632 VSS.n2631 0.0545365
R4420 VSS.n490 VSS.n482 0.0545365
R4421 VSS.n2327 VSS.n134 0.0545365
R4422 VSS.n1482 VSS.n651 0.048119
R4423 VSS.n1483 VSS.n1482 0.048119
R4424 VSS.n1401 VSS.n582 0.048119
R4425 VSS.n1393 VSS.n582 0.048119
R4426 VSS.n1077 VSS.n1076 0.048119
R4427 VSS.n1076 VSS.n881 0.048119
R4428 VSS.n2349 VSS.n127 0.048119
R4429 VSS.n2349 VSS.n2348 0.048119
R4430 VSS.n1083 VSS.n1082 0.048119
R4431 VSS.n1423 VSS.n696 0.048119
R4432 VSS.n2328 VSS.n133 0.0325513
R4433 VSS.n2642 VSS.n10 0.0281615
R4434 VSS.n492 VSS.n483 0.0281615
R4435 VSS.n2325 VSS.n135 0.0281615
R4436 VSS.n2345 VSS.n129 0.0265417
R4437 VSS.n2335 VSS.n129 0.0265417
R4438 VSS.n9 VSS.n8 0.0265417
R4439 VSS.n2637 VSS.n2636 0.0265417
R4440 VSS.n491 VSS.n489 0.0265417
R4441 VSS.n497 VSS.n480 0.0265417
R4442 VSS.n2321 VSS.n2320 0.0265417
R4443 VSS.n2326 VSS.n132 0.0265417
R4444 VSS.n3 VSS.n2 0.0265417
R4445 VSS.n4 VSS.n3 0.0265417
R4446 VSS.n2339 VSS.n2333 0.0257135
R4447 VSS.n2653 VSS.n5 0.0257135
R4448 VSS.n2632 VSS.n9 0.0200312
R4449 VSS.n491 VSS.n490 0.0200312
R4450 VSS.n2327 VSS.n2326 0.0200312
R4451 VSS.n8 VSS.n7 0.0174271
R4452 VSS.n2637 VSS.n13 0.0174271
R4453 VSS.n489 VSS.n488 0.0174271
R4454 VSS.n498 VSS.n497 0.0174271
R4455 VSS.n2320 VSS.n2319 0.0174271
R4456 VSS.n2329 VSS.n132 0.0174271
R4457 VSS.n2324 VSS.n2323 0.0165939
R4458 VSS.n2641 VSS.n2640 0.0165939
R4459 VSS.n494 VSS.n493 0.0165939
R4460 VSS.n2341 VSS.n2340 0.0151697
R4461 VSS.n2652 VSS.n2651 0.0151697
R4462 VSS.n2318 VSS.n133 0.0123942
R4463 VSS.n2635 VSS.n2634 0.010504
R4464 VSS.n2344 VSS.n2343 0.0102917
R4465 VSS.n2343 VSS.n2333 0.0102917
R4466 VSS.n2339 VSS.n2338 0.0102917
R4467 VSS.n2644 VSS.n2643 0.0102917
R4468 VSS.n2643 VSS.n2642 0.0102917
R4469 VSS.n2638 VSS.n10 0.0102917
R4470 VSS.n2638 VSS.n12 0.0102917
R4471 VSS.n487 VSS.n485 0.0102917
R4472 VSS.n492 VSS.n485 0.0102917
R4473 VSS.n496 VSS.n483 0.0102917
R4474 VSS.n136 VSS.n135 0.0102917
R4475 VSS.n2325 VSS.n131 0.0102917
R4476 VSS.n2330 VSS.n131 0.0102917
R4477 VSS.n2655 VSS.n2654 0.0102917
R4478 VSS.n2654 VSS.n2653 0.0102917
R4479 VSS.n2649 VSS.n5 0.0102917
R4480 VSS.n2631 VSS.n13 0.00961458
R4481 VSS.n498 VSS.n482 0.00961458
R4482 VSS.n2319 VSS.n134 0.00961458
R4483 VSS.n496 VSS.n495 0.00750807
R4484 VSS.n2322 VSS.n136 0.00750807
R4485 VSS.n2338 VSS.n2337 0.00748237
R4486 VSS.n2649 VSS.n2648 0.00748237
R4487 VSS.n2324 VSS.n130 0.00619697
R4488 VSS.n2331 VSS.n130 0.00619697
R4489 VSS.n2342 VSS.n2332 0.00619697
R4490 VSS.n2342 VSS.n2341 0.00619697
R4491 VSS.n2340 VSS.n2334 0.00619697
R4492 VSS.n2334 VSS.n0 0.00619697
R4493 VSS.n2656 VSS.n1 0.00619697
R4494 VSS.n2652 VSS.n1 0.00619697
R4495 VSS.n2651 VSS.n2650 0.00619697
R4496 VSS.n2650 VSS.n2646 0.00619697
R4497 VSS.n2645 VSS.n6 0.00619697
R4498 VSS.n2641 VSS.n6 0.00619697
R4499 VSS.n2640 VSS.n2639 0.00619697
R4500 VSS.n2639 VSS.n11 0.00619697
R4501 VSS.n486 VSS.n484 0.00619697
R4502 VSS.n493 VSS.n484 0.00619697
R4503 VSS.n2634 VSS.n2633 0.00370513
R4504 a_2479_7336.n0 a_2479_7336.t31 260.486
R4505 a_2479_7336.n68 a_2479_7336.t19 260.486
R4506 a_2479_7336.n79 a_2479_7336.t34 260.111
R4507 a_2479_7336.n80 a_2479_7336.t21 260.111
R4508 a_2479_7336.n81 a_2479_7336.t29 260.111
R4509 a_2479_7336.n82 a_2479_7336.t18 260.111
R4510 a_2479_7336.n83 a_2479_7336.t33 260.111
R4511 a_2479_7336.n84 a_2479_7336.t27 260.111
R4512 a_2479_7336.n1 a_2479_7336.t24 260.111
R4513 a_2479_7336.n0 a_2479_7336.t22 260.111
R4514 a_2479_7336.n68 a_2479_7336.t28 260.111
R4515 a_2479_7336.n69 a_2479_7336.t35 260.111
R4516 a_2479_7336.n71 a_2479_7336.t32 260.111
R4517 a_2479_7336.n72 a_2479_7336.t26 260.111
R4518 a_2479_7336.n73 a_2479_7336.t23 260.111
R4519 a_2479_7336.n74 a_2479_7336.t20 260.111
R4520 a_2479_7336.n75 a_2479_7336.t30 260.111
R4521 a_2479_7336.n76 a_2479_7336.t25 260.111
R4522 a_2479_7336.n86 a_2479_7336.n85 203.843
R4523 a_2479_7336.n70 a_2479_7336.n67 203.843
R4524 a_2479_7336.n59 a_2479_7336.n41 185
R4525 a_2479_7336.n59 a_2479_7336.n40 185
R4526 a_2479_7336.n59 a_2479_7336.n39 185
R4527 a_2479_7336.n59 a_2479_7336.n38 185
R4528 a_2479_7336.n59 a_2479_7336.n37 185
R4529 a_2479_7336.n59 a_2479_7336.n36 185
R4530 a_2479_7336.n59 a_2479_7336.n35 185
R4531 a_2479_7336.n28 a_2479_7336.n10 185
R4532 a_2479_7336.n28 a_2479_7336.n9 185
R4533 a_2479_7336.n28 a_2479_7336.n8 185
R4534 a_2479_7336.n28 a_2479_7336.n7 185
R4535 a_2479_7336.n28 a_2479_7336.n6 185
R4536 a_2479_7336.n28 a_2479_7336.n5 185
R4537 a_2479_7336.n28 a_2479_7336.n4 185
R4538 a_2479_7336.n43 a_2479_7336.t10 130.75
R4539 a_2479_7336.n12 a_2479_7336.t13 130.75
R4540 a_2479_7336.n43 a_2479_7336.t12 91.3557
R4541 a_2479_7336.n12 a_2479_7336.t14 91.3557
R4542 a_2479_7336.n60 a_2479_7336.n59 86.5152
R4543 a_2479_7336.n29 a_2479_7336.n28 86.5152
R4544 a_2479_7336.n58 a_2479_7336.n42 30.3012
R4545 a_2479_7336.n27 a_2479_7336.n11 30.3012
R4546 a_2479_7336.n67 a_2479_7336.t17 28.5655
R4547 a_2479_7336.n67 a_2479_7336.t1 28.5655
R4548 a_2479_7336.n86 a_2479_7336.t9 28.5655
R4549 a_2479_7336.t0 a_2479_7336.n86 28.5655
R4550 a_2479_7336.n35 a_2479_7336.n34 24.8476
R4551 a_2479_7336.n4 a_2479_7336.n3 24.8476
R4552 a_2479_7336.n44 a_2479_7336.n36 23.3417
R4553 a_2479_7336.n13 a_2479_7336.n5 23.3417
R4554 a_2479_7336.n61 a_2479_7336.n60 22.0256
R4555 a_2479_7336.n30 a_2479_7336.n29 22.0256
R4556 a_2479_7336.n46 a_2479_7336.n37 21.8358
R4557 a_2479_7336.n15 a_2479_7336.n6 21.8358
R4558 a_2479_7336.n48 a_2479_7336.n38 20.3299
R4559 a_2479_7336.n17 a_2479_7336.n7 20.3299
R4560 a_2479_7336.n50 a_2479_7336.n39 18.824
R4561 a_2479_7336.n19 a_2479_7336.n8 18.824
R4562 a_2479_7336.n52 a_2479_7336.n40 17.3181
R4563 a_2479_7336.n21 a_2479_7336.n9 17.3181
R4564 a_2479_7336.n59 a_2479_7336.n58 16.3559
R4565 a_2479_7336.n28 a_2479_7336.n27 16.3559
R4566 a_2479_7336.n54 a_2479_7336.n41 15.8123
R4567 a_2479_7336.n23 a_2479_7336.n10 15.8123
R4568 a_2479_7336.n64 a_2479_7336.n63 14.6052
R4569 a_2479_7336.n66 a_2479_7336.n65 14.6052
R4570 a_2479_7336.n32 a_2479_7336.n31 14.377
R4571 a_2479_7336.n60 a_2479_7336.n34 12.7256
R4572 a_2479_7336.n29 a_2479_7336.n3 12.7256
R4573 a_2479_7336.n77 a_2479_7336.t8 12.5928
R4574 a_2479_7336.n64 a_2479_7336.n62 11.5586
R4575 a_2479_7336.n42 a_2479_7336.n41 11.2946
R4576 a_2479_7336.n11 a_2479_7336.n10 11.2946
R4577 a_2479_7336.n54 a_2479_7336.n40 9.78874
R4578 a_2479_7336.n23 a_2479_7336.n9 9.78874
R4579 a_2479_7336.n34 a_2479_7336.n33 9.3005
R4580 a_2479_7336.n45 a_2479_7336.n44 9.3005
R4581 a_2479_7336.n47 a_2479_7336.n46 9.3005
R4582 a_2479_7336.n49 a_2479_7336.n48 9.3005
R4583 a_2479_7336.n51 a_2479_7336.n50 9.3005
R4584 a_2479_7336.n53 a_2479_7336.n52 9.3005
R4585 a_2479_7336.n55 a_2479_7336.n54 9.3005
R4586 a_2479_7336.n56 a_2479_7336.n42 9.3005
R4587 a_2479_7336.n3 a_2479_7336.n2 9.3005
R4588 a_2479_7336.n14 a_2479_7336.n13 9.3005
R4589 a_2479_7336.n16 a_2479_7336.n15 9.3005
R4590 a_2479_7336.n18 a_2479_7336.n17 9.3005
R4591 a_2479_7336.n20 a_2479_7336.n19 9.3005
R4592 a_2479_7336.n22 a_2479_7336.n21 9.3005
R4593 a_2479_7336.n24 a_2479_7336.n23 9.3005
R4594 a_2479_7336.n25 a_2479_7336.n11 9.3005
R4595 a_2479_7336.n52 a_2479_7336.n39 8.28285
R4596 a_2479_7336.n21 a_2479_7336.n8 8.28285
R4597 a_2479_7336.n78 a_2479_7336.n66 7.17277
R4598 a_2479_7336.n50 a_2479_7336.n38 6.77697
R4599 a_2479_7336.n19 a_2479_7336.n7 6.77697
R4600 a_2479_7336.n32 a_2479_7336.n30 6.19091
R4601 a_2479_7336.n48 a_2479_7336.n37 5.27109
R4602 a_2479_7336.n17 a_2479_7336.n6 5.27109
R4603 a_2479_7336.n78 a_2479_7336.n77 4.74179
R4604 a_2479_7336.n46 a_2479_7336.n36 3.76521
R4605 a_2479_7336.n15 a_2479_7336.n5 3.76521
R4606 a_2479_7336.n62 a_2479_7336.n61 3.31388
R4607 a_2479_7336.n66 a_2479_7336.n64 2.87753
R4608 a_2479_7336.n63 a_2479_7336.t5 2.48621
R4609 a_2479_7336.n63 a_2479_7336.t4 2.48621
R4610 a_2479_7336.n65 a_2479_7336.t3 2.48621
R4611 a_2479_7336.n65 a_2479_7336.t2 2.48621
R4612 a_2479_7336.n59 a_2479_7336.t15 2.48621
R4613 a_2479_7336.n59 a_2479_7336.t11 2.48621
R4614 a_2479_7336.n28 a_2479_7336.t14 2.48621
R4615 a_2479_7336.n28 a_2479_7336.t7 2.48621
R4616 a_2479_7336.n31 a_2479_7336.t16 2.48621
R4617 a_2479_7336.n31 a_2479_7336.t6 2.48621
R4618 a_2479_7336.n58 a_2479_7336.n57 2.36936
R4619 a_2479_7336.n27 a_2479_7336.n26 2.36936
R4620 a_2479_7336.n62 a_2479_7336.n32 2.30287
R4621 a_2479_7336.n44 a_2479_7336.n35 2.25932
R4622 a_2479_7336.n13 a_2479_7336.n4 2.25932
R4623 a_2479_7336.n77 a_2479_7336.n76 1.41083
R4624 a_2479_7336.n79 a_2479_7336.n78 1.23683
R4625 a_2479_7336.n76 a_2479_7336.n75 0.3755
R4626 a_2479_7336.n75 a_2479_7336.n74 0.3755
R4627 a_2479_7336.n74 a_2479_7336.n73 0.3755
R4628 a_2479_7336.n73 a_2479_7336.n72 0.3755
R4629 a_2479_7336.n72 a_2479_7336.n71 0.3755
R4630 a_2479_7336.n69 a_2479_7336.n68 0.3755
R4631 a_2479_7336.n1 a_2479_7336.n0 0.3755
R4632 a_2479_7336.n84 a_2479_7336.n83 0.3755
R4633 a_2479_7336.n83 a_2479_7336.n82 0.3755
R4634 a_2479_7336.n82 a_2479_7336.n81 0.3755
R4635 a_2479_7336.n81 a_2479_7336.n80 0.3755
R4636 a_2479_7336.n80 a_2479_7336.n79 0.3755
R4637 a_2479_7336.n57 a_2479_7336.n43 0.320353
R4638 a_2479_7336.n26 a_2479_7336.n12 0.320353
R4639 a_2479_7336.n57 a_2479_7336.n56 0.196152
R4640 a_2479_7336.n56 a_2479_7336.n55 0.196152
R4641 a_2479_7336.n55 a_2479_7336.n53 0.196152
R4642 a_2479_7336.n53 a_2479_7336.n51 0.196152
R4643 a_2479_7336.n51 a_2479_7336.n49 0.196152
R4644 a_2479_7336.n49 a_2479_7336.n47 0.196152
R4645 a_2479_7336.n47 a_2479_7336.n45 0.196152
R4646 a_2479_7336.n45 a_2479_7336.n33 0.196152
R4647 a_2479_7336.n61 a_2479_7336.n33 0.196152
R4648 a_2479_7336.n26 a_2479_7336.n25 0.196152
R4649 a_2479_7336.n25 a_2479_7336.n24 0.196152
R4650 a_2479_7336.n24 a_2479_7336.n22 0.196152
R4651 a_2479_7336.n22 a_2479_7336.n20 0.196152
R4652 a_2479_7336.n20 a_2479_7336.n18 0.196152
R4653 a_2479_7336.n18 a_2479_7336.n16 0.196152
R4654 a_2479_7336.n16 a_2479_7336.n14 0.196152
R4655 a_2479_7336.n14 a_2479_7336.n2 0.196152
R4656 a_2479_7336.n30 a_2479_7336.n2 0.196152
R4657 a_2479_7336.n71 a_2479_7336.n70 0.188
R4658 a_2479_7336.n70 a_2479_7336.n69 0.188
R4659 a_2479_7336.n85 a_2479_7336.n1 0.188
R4660 a_2479_7336.n85 a_2479_7336.n84 0.188
R4661 VOUT.n13 VOUT.t8 260.298
R4662 VOUT.t4 VOUT.n13 260.298
R4663 VOUT.t8 VOUT.n8 260.298
R4664 VOUT.n56 VOUT.t6 260.298
R4665 VOUT.t2 VOUT.n56 260.298
R4666 VOUT.n57 VOUT.t2 260.298
R4667 VOUT.n14 VOUT.t4 260.111
R4668 VOUT.t6 VOUT.n54 260.111
R4669 VOUT.n12 VOUT.t10 232.03
R4670 VOUT.t3 VOUT.n55 232.03
R4671 VOUT.n2 VOUT.n0 206.708
R4672 VOUT.n6 VOUT.n5 206.094
R4673 VOUT.n4 VOUT.n3 206.094
R4674 VOUT.n2 VOUT.n1 206.094
R4675 VOUT.n70 VOUT.n69 206.094
R4676 VOUT.n68 VOUT.n67 206.094
R4677 VOUT.n66 VOUT.n65 206.094
R4678 VOUT.n64 VOUT.n63 206.094
R4679 VOUT.n11 VOUT.n10 203.03
R4680 VOUT.n9 VOUT.n7 203.03
R4681 VOUT.n61 VOUT.n60 203.03
R4682 VOUT.n59 VOUT.n58 203.03
R4683 VOUT.n43 VOUT.n42 185
R4684 VOUT.n43 VOUT.n25 185
R4685 VOUT.n43 VOUT.n24 185
R4686 VOUT.n43 VOUT.n23 185
R4687 VOUT.n43 VOUT.n22 185
R4688 VOUT.n43 VOUT.n21 185
R4689 VOUT.n43 VOUT.n20 185
R4690 VOUT.n26 VOUT.t11 130.75
R4691 VOUT.n26 VOUT.t13 91.3557
R4692 VOUT.n44 VOUT.n43 86.5152
R4693 VOUT.n28 VOUT.n19 30.3012
R4694 VOUT.n10 VOUT.t5 28.5655
R4695 VOUT.n10 VOUT.t9 28.5655
R4696 VOUT.n9 VOUT.t24 28.5655
R4697 VOUT.t5 VOUT.n9 28.5655
R4698 VOUT.n5 VOUT.t21 28.5655
R4699 VOUT.n5 VOUT.t30 28.5655
R4700 VOUT.n3 VOUT.t23 28.5655
R4701 VOUT.n3 VOUT.t31 28.5655
R4702 VOUT.n1 VOUT.t25 28.5655
R4703 VOUT.n1 VOUT.t14 28.5655
R4704 VOUT.n0 VOUT.t27 28.5655
R4705 VOUT.n0 VOUT.t28 28.5655
R4706 VOUT.n60 VOUT.t7 28.5655
R4707 VOUT.n60 VOUT.t17 28.5655
R4708 VOUT.n59 VOUT.t3 28.5655
R4709 VOUT.t7 VOUT.n59 28.5655
R4710 VOUT.n69 VOUT.t18 28.5655
R4711 VOUT.n69 VOUT.t20 28.5655
R4712 VOUT.n67 VOUT.t26 28.5655
R4713 VOUT.n67 VOUT.t29 28.5655
R4714 VOUT.n65 VOUT.t22 28.5655
R4715 VOUT.n65 VOUT.t19 28.5655
R4716 VOUT.n63 VOUT.t15 28.5655
R4717 VOUT.n63 VOUT.t16 28.5655
R4718 VOUT.n42 VOUT.n18 24.8476
R4719 VOUT.n41 VOUT.n25 23.3417
R4720 VOUT.n45 VOUT.n44 22.0256
R4721 VOUT.n38 VOUT.n24 21.8358
R4722 VOUT.n36 VOUT.n23 20.3299
R4723 VOUT.n46 VOUT.n45 19.0885
R4724 VOUT.n34 VOUT.n22 18.824
R4725 VOUT.n32 VOUT.n21 17.3181
R4726 VOUT.n43 VOUT.n19 16.3559
R4727 VOUT.n30 VOUT.n20 15.8123
R4728 VOUT.n44 VOUT.n18 12.7256
R4729 VOUT.n28 VOUT.n20 11.2946
R4730 VOUT.n30 VOUT.n21 9.78874
R4731 VOUT.n18 VOUT.n17 9.3005
R4732 VOUT.n41 VOUT.n40 9.3005
R4733 VOUT.n39 VOUT.n38 9.3005
R4734 VOUT.n37 VOUT.n36 9.3005
R4735 VOUT.n35 VOUT.n34 9.3005
R4736 VOUT.n33 VOUT.n32 9.3005
R4737 VOUT.n31 VOUT.n30 9.3005
R4738 VOUT.n29 VOUT.n28 9.3005
R4739 VOUT.n32 VOUT.n22 8.28285
R4740 VOUT.n34 VOUT.n23 6.77697
R4741 VOUT.n36 VOUT.n24 5.27109
R4742 VOUT.n38 VOUT.n25 3.76521
R4743 VOUT.n48 VOUT.n47 3.4105
R4744 VOUT.n72 VOUT.n46 3.29996
R4745 VOUT.n64 VOUT.n62 3.23261
R4746 VOUT.n16 VOUT.n15 2.55612
R4747 VOUT.n43 VOUT.t0 2.48621
R4748 VOUT.n43 VOUT.t12 2.48621
R4749 VOUT VOUT.n16 2.47337
R4750 VOUT.n27 VOUT.n19 2.36936
R4751 VOUT.n42 VOUT.n41 2.25932
R4752 VOUT.n71 VOUT.n70 2.12962
R4753 VOUT.n53 VOUT.n52 1.70927
R4754 VOUT.n51 VOUT.n50 1.7055
R4755 VOUT.n50 VOUT.n49 1.7055
R4756 VOUT.n52 VOUT.n51 1.14963
R4757 VOUT.n72 VOUT.n71 1.09816
R4758 VOUT.n4 VOUT.n2 0.61449
R4759 VOUT.n6 VOUT.n4 0.61449
R4760 VOUT.n16 VOUT.n6 0.61449
R4761 VOUT.n66 VOUT.n64 0.61449
R4762 VOUT.n68 VOUT.n66 0.61449
R4763 VOUT.n70 VOUT.n68 0.61449
R4764 VOUT.n51 VOUT.t1 0.563396
R4765 VOUT VOUT.n72 0.521984
R4766 VOUT.n62 VOUT.n61 0.446229
R4767 VOUT.n61 VOUT.n55 0.43664
R4768 VOUT.n12 VOUT.n7 0.436638
R4769 VOUT.n15 VOUT.n7 0.38373
R4770 VOUT.n11 VOUT.n8 0.38373
R4771 VOUT.n58 VOUT.n57 0.383729
R4772 VOUT.n27 VOUT.n26 0.320353
R4773 VOUT.n13 VOUT.n12 0.285826
R4774 VOUT.n56 VOUT.n55 0.285826
R4775 VOUT.n49 VOUT.n46 0.2193
R4776 VOUT.n45 VOUT.n17 0.196152
R4777 VOUT.n40 VOUT.n17 0.196152
R4778 VOUT.n40 VOUT.n39 0.196152
R4779 VOUT.n39 VOUT.n37 0.196152
R4780 VOUT.n37 VOUT.n35 0.196152
R4781 VOUT.n35 VOUT.n33 0.196152
R4782 VOUT.n33 VOUT.n31 0.196152
R4783 VOUT.n31 VOUT.n29 0.196152
R4784 VOUT.n29 VOUT.n27 0.196152
R4785 VOUT.n15 VOUT.n14 0.188
R4786 VOUT.n14 VOUT.n8 0.188
R4787 VOUT.n57 VOUT.n54 0.188
R4788 VOUT.n62 VOUT.n54 0.1255
R4789 VOUT.n58 VOUT.n55 0.0984044
R4790 VOUT.n12 VOUT.n11 0.0984028
R4791 VOUT.n71 VOUT.n53 0.0647077
R4792 VOUT.n50 VOUT.n48 0.0102917
R4793 VOUT.n52 VOUT.n48 0.00750288
R4794 VOUT.n53 VOUT.n47 0.00118306
R4795 VOUT.n49 VOUT.n47 0.00118306
R4796 VDD.n256 VDD.n153 723.529
R4797 VDD.n168 VDD.n156 723.529
R4798 VDD.n311 VDD.n19 723.529
R4799 VDD.n115 VDD.n24 723.529
R4800 VDD.n230 VDD.n229 515.294
R4801 VDD.n245 VDD.n244 275.295
R4802 VDD.n321 VDD.n14 275.295
R4803 VDD.n350 VDD.t16 260.486
R4804 VDD.n334 VDD.t36 260.486
R4805 VDD.n39 VDD.t52 260.486
R4806 VDD.n64 VDD.t27 260.486
R4807 VDD.t22 VDD.n347 260.298
R4808 VDD.t40 VDD.n349 260.298
R4809 VDD.n354 VDD.t22 260.298
R4810 VDD.n331 VDD.t47 260.298
R4811 VDD.t47 VDD.n328 260.298
R4812 VDD.n335 VDD.t54 260.298
R4813 VDD.t9 VDD.n43 260.298
R4814 VDD.n41 VDD.t30 260.298
R4815 VDD.n44 VDD.t9 260.298
R4816 VDD.t49 VDD.n63 260.298
R4817 VDD.n61 VDD.t38 260.298
R4818 VDD.n57 VDD.t38 260.298
R4819 VDD.n1 VDD.t19 260.199
R4820 VDD.n372 VDD.t42 260.199
R4821 VDD.n353 VDD.t45 260.111
R4822 VDD.t45 VDD.n352 260.111
R4823 VDD.n350 VDD.t40 260.111
R4824 VDD.t54 VDD.n334 260.111
R4825 VDD.n333 VDD.t25 260.111
R4826 VDD.t25 VDD.n332 260.111
R4827 VDD.t33 VDD.n37 260.111
R4828 VDD.n42 VDD.t33 260.111
R4829 VDD.t30 VDD.n39 260.111
R4830 VDD.n64 VDD.t49 260.111
R4831 VDD.t13 VDD.n56 260.111
R4832 VDD.n62 VDD.t13 260.111
R4833 VDD.n170 VDD.n169 240
R4834 VDD.n173 VDD.n169 240
R4835 VDD.n249 VDD.n248 240
R4836 VDD.n237 VDD.n236 240
R4837 VDD.n234 VDD.n233 240
R4838 VDD.n226 VDD.n225 240
R4839 VDD.n222 VDD.n221 240
R4840 VDD.n218 VDD.n217 240
R4841 VDD.n214 VDD.n213 240
R4842 VDD.n210 VDD.n209 240
R4843 VDD.n206 VDD.n168 240
R4844 VDD.n307 VDD.n19 240
R4845 VDD.n307 VDD.n21 240
R4846 VDD.n120 VDD.n21 240
R4847 VDD.n121 VDD.n120 240
R4848 VDD.n122 VDD.n121 240
R4849 VDD.n181 VDD.n122 240
R4850 VDD.n181 VDD.n127 240
R4851 VDD.n128 VDD.n127 240
R4852 VDD.n129 VDD.n128 240
R4853 VDD.n186 VDD.n129 240
R4854 VDD.n186 VDD.n134 240
R4855 VDD.n135 VDD.n134 240
R4856 VDD.n136 VDD.n135 240
R4857 VDD.n191 VDD.n136 240
R4858 VDD.n191 VDD.n141 240
R4859 VDD.n142 VDD.n141 240
R4860 VDD.n143 VDD.n142 240
R4861 VDD.n196 VDD.n143 240
R4862 VDD.n196 VDD.n148 240
R4863 VDD.n149 VDD.n148 240
R4864 VDD.n150 VDD.n149 240
R4865 VDD.n201 VDD.n150 240
R4866 VDD.n201 VDD.n155 240
R4867 VDD.n156 VDD.n155 240
R4868 VDD.n113 VDD.n112 240
R4869 VDD.n110 VDD.n28 240
R4870 VDD.n106 VDD.n105 240
R4871 VDD.n103 VDD.n31 240
R4872 VDD.n97 VDD.n96 240
R4873 VDD.n94 VDD.n75 240
R4874 VDD.n90 VDD.n89 240
R4875 VDD.n87 VDD.n78 240
R4876 VDD.n83 VDD.n82 240
R4877 VDD.n319 VDD.n16 240
R4878 VDD.n314 VDD.n313 240
R4879 VDD.n305 VDD.n24 240
R4880 VDD.n305 VDD.n25 240
R4881 VDD.n301 VDD.n25 240
R4882 VDD.n301 VDD.n119 240
R4883 VDD.n297 VDD.n119 240
R4884 VDD.n297 VDD.n124 240
R4885 VDD.n293 VDD.n124 240
R4886 VDD.n293 VDD.n126 240
R4887 VDD.n289 VDD.n126 240
R4888 VDD.n289 VDD.n131 240
R4889 VDD.n285 VDD.n131 240
R4890 VDD.n285 VDD.n133 240
R4891 VDD.n281 VDD.n133 240
R4892 VDD.n281 VDD.n137 240
R4893 VDD.n277 VDD.n137 240
R4894 VDD.n277 VDD.n139 240
R4895 VDD.n273 VDD.n139 240
R4896 VDD.n273 VDD.n144 240
R4897 VDD.n269 VDD.n144 240
R4898 VDD.n269 VDD.n146 240
R4899 VDD.n265 VDD.n146 240
R4900 VDD.n265 VDD.n151 240
R4901 VDD.n261 VDD.n151 240
R4902 VDD.n261 VDD.n153 240
R4903 VDD.n355 VDD.t24 232.03
R4904 VDD.t48 VDD.n327 232.03
R4905 VDD.n36 VDD.t12 232.03
R4906 VDD.n60 VDD.t39 232.03
R4907 VDD.n371 VDD.t44 231.758
R4908 VDD.n365 VDD.n363 206.48
R4909 VDD.n344 VDD.n343 205.865
R4910 VDD.n369 VDD.n368 205.865
R4911 VDD.n367 VDD.n366 205.865
R4912 VDD.n365 VDD.n364 205.865
R4913 VDD.n9 VDD.n8 205.865
R4914 VDD.n7 VDD.n6 205.865
R4915 VDD.n5 VDD.n4 205.865
R4916 VDD.n3 VDD.n2 205.865
R4917 VDD.n53 VDD.n52 205.865
R4918 VDD.n371 VDD.n370 203.143
R4919 VDD.n361 VDD.n360 203.127
R4920 VDD.n341 VDD.n340 203.127
R4921 VDD.n50 VDD.n49 203.127
R4922 VDD.n70 VDD.n69 203.127
R4923 VDD.n359 VDD.n345 203.126
R4924 VDD.n339 VDD.n325 203.126
R4925 VDD.n48 VDD.n34 203.126
R4926 VDD.n68 VDD.n54 203.126
R4927 VDD.n358 VDD.n346 203.03
R4928 VDD.n357 VDD.n356 203.03
R4929 VDD.n338 VDD.n337 203.03
R4930 VDD.n330 VDD.n329 203.03
R4931 VDD.n47 VDD.n35 203.03
R4932 VDD.n46 VDD.n45 203.03
R4933 VDD.n67 VDD.n66 203.03
R4934 VDD.n59 VDD.n58 203.03
R4935 VDD.n117 VDD.n24 185
R4936 VDD.n24 VDD.n23 185
R4937 VDD.n305 VDD.n304 185
R4938 VDD.n306 VDD.n305 185
R4939 VDD.n303 VDD.n25 185
R4940 VDD.n25 VDD.n22 185
R4941 VDD.n302 VDD.n301 185
R4942 VDD.n301 VDD.n300 185
R4943 VDD.n119 VDD.n118 185
R4944 VDD.n299 VDD.n119 185
R4945 VDD.n297 VDD.n296 185
R4946 VDD.n298 VDD.n297 185
R4947 VDD.n295 VDD.n124 185
R4948 VDD.n124 VDD.n123 185
R4949 VDD.n294 VDD.n293 185
R4950 VDD.n293 VDD.n292 185
R4951 VDD.n126 VDD.n125 185
R4952 VDD.n291 VDD.n126 185
R4953 VDD.n289 VDD.n288 185
R4954 VDD.n290 VDD.n289 185
R4955 VDD.n287 VDD.n131 185
R4956 VDD.n131 VDD.n130 185
R4957 VDD.n286 VDD.n285 185
R4958 VDD.n285 VDD.n284 185
R4959 VDD.n133 VDD.n132 185
R4960 VDD.n283 VDD.n133 185
R4961 VDD.n281 VDD.n280 185
R4962 VDD.n282 VDD.n281 185
R4963 VDD.n279 VDD.n137 185
R4964 VDD.n140 VDD.n137 185
R4965 VDD.n278 VDD.n277 185
R4966 VDD.n277 VDD.n276 185
R4967 VDD.n139 VDD.n138 185
R4968 VDD.n275 VDD.n139 185
R4969 VDD.n273 VDD.n272 185
R4970 VDD.n274 VDD.n273 185
R4971 VDD.n271 VDD.n144 185
R4972 VDD.n147 VDD.n144 185
R4973 VDD.n270 VDD.n269 185
R4974 VDD.n269 VDD.n268 185
R4975 VDD.n146 VDD.n145 185
R4976 VDD.n267 VDD.n146 185
R4977 VDD.n265 VDD.n264 185
R4978 VDD.n266 VDD.n265 185
R4979 VDD.n263 VDD.n151 185
R4980 VDD.n154 VDD.n151 185
R4981 VDD.n262 VDD.n261 185
R4982 VDD.n261 VDD.n260 185
R4983 VDD.n153 VDD.n152 185
R4984 VDD.n259 VDD.n153 185
R4985 VDD.n256 VDD.n255 185
R4986 VDD.n254 VDD.n170 185
R4987 VDD.n171 VDD.n169 185
R4988 VDD.n258 VDD.n169 185
R4989 VDD.n174 VDD.n173 185
R4990 VDD.n250 VDD.n249 185
R4991 VDD.n248 VDD.n247 185
R4992 VDD.n246 VDD.n245 185
R4993 VDD.n244 VDD.n243 185
R4994 VDD.n236 VDD.n175 185
R4995 VDD.n238 VDD.n237 185
R4996 VDD.n235 VDD.n234 185
R4997 VDD.n233 VDD.n232 185
R4998 VDD.n231 VDD.n230 185
R4999 VDD.n229 VDD.n228 185
R5000 VDD.n227 VDD.n226 185
R5001 VDD.n225 VDD.n224 185
R5002 VDD.n223 VDD.n222 185
R5003 VDD.n221 VDD.n220 185
R5004 VDD.n219 VDD.n218 185
R5005 VDD.n217 VDD.n216 185
R5006 VDD.n215 VDD.n214 185
R5007 VDD.n213 VDD.n212 185
R5008 VDD.n211 VDD.n210 185
R5009 VDD.n209 VDD.n208 185
R5010 VDD.n207 VDD.n206 185
R5011 VDD.n205 VDD.n168 185
R5012 VDD.n258 VDD.n168 185
R5013 VDD.n204 VDD.n156 185
R5014 VDD.n259 VDD.n156 185
R5015 VDD.n203 VDD.n155 185
R5016 VDD.n260 VDD.n155 185
R5017 VDD.n202 VDD.n201 185
R5018 VDD.n201 VDD.n154 185
R5019 VDD.n200 VDD.n150 185
R5020 VDD.n266 VDD.n150 185
R5021 VDD.n199 VDD.n149 185
R5022 VDD.n267 VDD.n149 185
R5023 VDD.n198 VDD.n148 185
R5024 VDD.n268 VDD.n148 185
R5025 VDD.n197 VDD.n196 185
R5026 VDD.n196 VDD.n147 185
R5027 VDD.n195 VDD.n143 185
R5028 VDD.n274 VDD.n143 185
R5029 VDD.n194 VDD.n142 185
R5030 VDD.n275 VDD.n142 185
R5031 VDD.n193 VDD.n141 185
R5032 VDD.n276 VDD.n141 185
R5033 VDD.n192 VDD.n191 185
R5034 VDD.n191 VDD.n140 185
R5035 VDD.n190 VDD.n136 185
R5036 VDD.n282 VDD.n136 185
R5037 VDD.n189 VDD.n135 185
R5038 VDD.n283 VDD.n135 185
R5039 VDD.n188 VDD.n134 185
R5040 VDD.n284 VDD.n134 185
R5041 VDD.n187 VDD.n186 185
R5042 VDD.n186 VDD.n130 185
R5043 VDD.n185 VDD.n129 185
R5044 VDD.n290 VDD.n129 185
R5045 VDD.n184 VDD.n128 185
R5046 VDD.n291 VDD.n128 185
R5047 VDD.n183 VDD.n127 185
R5048 VDD.n292 VDD.n127 185
R5049 VDD.n182 VDD.n181 185
R5050 VDD.n181 VDD.n123 185
R5051 VDD.n180 VDD.n122 185
R5052 VDD.n298 VDD.n122 185
R5053 VDD.n179 VDD.n121 185
R5054 VDD.n299 VDD.n121 185
R5055 VDD.n178 VDD.n120 185
R5056 VDD.n300 VDD.n120 185
R5057 VDD.n21 VDD.n20 185
R5058 VDD.n22 VDD.n21 185
R5059 VDD.n308 VDD.n307 185
R5060 VDD.n307 VDD.n306 185
R5061 VDD.n309 VDD.n19 185
R5062 VDD.n23 VDD.n19 185
R5063 VDD.n311 VDD.n310 185
R5064 VDD.n313 VDD.n17 185
R5065 VDD.n315 VDD.n314 185
R5066 VDD.n316 VDD.n16 185
R5067 VDD.n319 VDD.n318 185
R5068 VDD.n322 VDD.n321 185
R5069 VDD.n14 VDD.n12 185
R5070 VDD.n82 VDD.n79 185
R5071 VDD.n84 VDD.n83 185
R5072 VDD.n85 VDD.n78 185
R5073 VDD.n87 VDD.n86 185
R5074 VDD.n89 VDD.n76 185
R5075 VDD.n91 VDD.n90 185
R5076 VDD.n92 VDD.n75 185
R5077 VDD.n94 VDD.n93 185
R5078 VDD.n96 VDD.n73 185
R5079 VDD.n98 VDD.n97 185
R5080 VDD.n33 VDD.n31 185
R5081 VDD.n103 VDD.n102 185
R5082 VDD.n105 VDD.n29 185
R5083 VDD.n107 VDD.n106 185
R5084 VDD.n108 VDD.n28 185
R5085 VDD.n110 VDD.n109 185
R5086 VDD.n112 VDD.n27 185
R5087 VDD.n113 VDD.n26 185
R5088 VDD.n116 VDD.n115 185
R5089 VDD.n90 VDD.n77 107.683
R5090 VDD.n77 VDD.n75 107.683
R5091 VDD.n1 VDD.n0 101.662
R5092 VDD.n217 VDD.n165 78.9253
R5093 VDD.n104 VDD.n103 78.9253
R5094 VDD.n214 VDD.n165 78.9253
R5095 VDD.n105 VDD.n104 78.9253
R5096 VDD.n117 VDD.n116 77.177
R5097 VDD.n255 VDD.n152 77.177
R5098 VDD.n205 VDD.n204 77.177
R5099 VDD.n310 VDD.n309 77.177
R5100 VDD.n257 VDD.n256 72.7879
R5101 VDD.n173 VDD.n157 72.7879
R5102 VDD.n248 VDD.n158 72.7879
R5103 VDD.n244 VDD.n159 72.7879
R5104 VDD.n237 VDD.n160 72.7879
R5105 VDD.n233 VDD.n161 72.7879
R5106 VDD.n229 VDD.n162 72.7879
R5107 VDD.n225 VDD.n163 72.7879
R5108 VDD.n221 VDD.n164 72.7879
R5109 VDD.n213 VDD.n166 72.7879
R5110 VDD.n209 VDD.n167 72.7879
R5111 VDD.n114 VDD.n113 72.7879
R5112 VDD.n111 VDD.n110 72.7879
R5113 VDD.n106 VDD.n30 72.7879
R5114 VDD.n97 VDD.n74 72.7879
R5115 VDD.n95 VDD.n94 72.7879
R5116 VDD.n88 VDD.n87 72.7879
R5117 VDD.n83 VDD.n80 72.7879
R5118 VDD.n81 VDD.n14 72.7879
R5119 VDD.n320 VDD.n319 72.7879
R5120 VDD.n314 VDD.n18 72.7879
R5121 VDD.n312 VDD.n311 72.7879
R5122 VDD.n257 VDD.n170 72.7879
R5123 VDD.n249 VDD.n157 72.7879
R5124 VDD.n245 VDD.n158 72.7879
R5125 VDD.n236 VDD.n159 72.7879
R5126 VDD.n234 VDD.n160 72.7879
R5127 VDD.n230 VDD.n161 72.7879
R5128 VDD.n226 VDD.n162 72.7879
R5129 VDD.n222 VDD.n163 72.7879
R5130 VDD.n218 VDD.n164 72.7879
R5131 VDD.n210 VDD.n166 72.7879
R5132 VDD.n206 VDD.n167 72.7879
R5133 VDD.n313 VDD.n312 72.7879
R5134 VDD.n18 VDD.n16 72.7879
R5135 VDD.n321 VDD.n320 72.7879
R5136 VDD.n82 VDD.n81 72.7879
R5137 VDD.n80 VDD.n78 72.7879
R5138 VDD.n89 VDD.n88 72.7879
R5139 VDD.n96 VDD.n95 72.7879
R5140 VDD.n74 VDD.n31 72.7879
R5141 VDD.n30 VDD.n28 72.7879
R5142 VDD.n112 VDD.n111 72.7879
R5143 VDD.n115 VDD.n114 72.7879
R5144 VDD.n23 VDD.n15 57.1093
R5145 VDD.n259 VDD.n258 57.1093
R5146 VDD.n258 VDD.n257 56.1076
R5147 VDD.n258 VDD.n157 56.1076
R5148 VDD.n258 VDD.n158 56.1076
R5149 VDD.n258 VDD.n159 56.1076
R5150 VDD.n258 VDD.n160 56.1076
R5151 VDD.n258 VDD.n161 56.1076
R5152 VDD.n258 VDD.n162 56.1076
R5153 VDD.n258 VDD.n163 56.1076
R5154 VDD.n258 VDD.n164 56.1076
R5155 VDD.n258 VDD.n166 56.1076
R5156 VDD.n258 VDD.n167 56.1076
R5157 VDD.n312 VDD.n15 56.1076
R5158 VDD.n18 VDD.n15 56.1076
R5159 VDD.n320 VDD.n15 56.1076
R5160 VDD.n81 VDD.n15 56.1076
R5161 VDD.n80 VDD.n15 56.1076
R5162 VDD.n88 VDD.n15 56.1076
R5163 VDD.n95 VDD.n15 56.1076
R5164 VDD.n74 VDD.n15 56.1076
R5165 VDD.n30 VDD.n15 56.1076
R5166 VDD.n111 VDD.n15 56.1076
R5167 VDD.n114 VDD.n15 56.1076
R5168 VDD.n231 VDD.n228 54.9652
R5169 VDD.n92 VDD.n91 54.9652
R5170 VDD.n258 VDD.n165 53.0388
R5171 VDD.n104 VDD.n15 53.0388
R5172 VDD.n0 VDD.t67 41.0864
R5173 VDD.n77 VDD.n15 38.6605
R5174 VDD.n306 VDD.n22 30.8211
R5175 VDD.n300 VDD.n299 30.8211
R5176 VDD.n298 VDD.n123 30.8211
R5177 VDD.n292 VDD.n291 30.8211
R5178 VDD.n290 VDD.n130 30.8211
R5179 VDD.n284 VDD.n283 30.8211
R5180 VDD.n283 VDD.n282 30.8211
R5181 VDD.n276 VDD.n140 30.8211
R5182 VDD.n275 VDD.n274 30.8211
R5183 VDD.n268 VDD.n147 30.8211
R5184 VDD.n267 VDD.n266 30.8211
R5185 VDD.n260 VDD.n154 30.8211
R5186 VDD.t0 VDD.n130 30.3679
R5187 VDD.n140 VDD.t7 30.3679
R5188 VDD.n291 VDD.t5 29.4614
R5189 VDD.t2 VDD.n275 29.4614
R5190 VDD.n246 VDD.n243 29.3652
R5191 VDD.n216 VDD.n215 29.3652
R5192 VDD.n8 VDD.t64 28.5655
R5193 VDD.n8 VDD.t73 28.5655
R5194 VDD.n6 VDD.t60 28.5655
R5195 VDD.n6 VDD.t57 28.5655
R5196 VDD.n4 VDD.t69 28.5655
R5197 VDD.n4 VDD.t66 28.5655
R5198 VDD.n2 VDD.t62 28.5655
R5199 VDD.n2 VDD.t72 28.5655
R5200 VDD.n360 VDD.t3 28.5655
R5201 VDD.n360 VDD.t18 28.5655
R5202 VDD.t41 VDD.n358 28.5655
R5203 VDD.n358 VDD.t46 28.5655
R5204 VDD.t46 VDD.n357 28.5655
R5205 VDD.n357 VDD.t23 28.5655
R5206 VDD.t18 VDD.n359 28.5655
R5207 VDD.n359 VDD.t41 28.5655
R5208 VDD.n340 VDD.t37 28.5655
R5209 VDD.n340 VDD.t56 28.5655
R5210 VDD.n338 VDD.t26 28.5655
R5211 VDD.t55 VDD.n338 28.5655
R5212 VDD.n329 VDD.t48 28.5655
R5213 VDD.n329 VDD.t26 28.5655
R5214 VDD.n339 VDD.t55 28.5655
R5215 VDD.t37 VDD.n339 28.5655
R5216 VDD.n343 VDD.t1 28.5655
R5217 VDD.n343 VDD.t8 28.5655
R5218 VDD.t32 VDD.n47 28.5655
R5219 VDD.n47 VDD.t35 28.5655
R5220 VDD.t35 VDD.n46 28.5655
R5221 VDD.n46 VDD.t11 28.5655
R5222 VDD.t53 VDD.n48 28.5655
R5223 VDD.n48 VDD.t32 28.5655
R5224 VDD.n49 VDD.t4 28.5655
R5225 VDD.n49 VDD.t53 28.5655
R5226 VDD.n52 VDD.t75 28.5655
R5227 VDD.n52 VDD.t76 28.5655
R5228 VDD.n67 VDD.t15 28.5655
R5229 VDD.t51 VDD.n67 28.5655
R5230 VDD.n58 VDD.t39 28.5655
R5231 VDD.n58 VDD.t15 28.5655
R5232 VDD.n68 VDD.t51 28.5655
R5233 VDD.t29 VDD.n68 28.5655
R5234 VDD.n69 VDD.t29 28.5655
R5235 VDD.n69 VDD.t6 28.5655
R5236 VDD.n370 VDD.t58 28.5655
R5237 VDD.n370 VDD.t43 28.5655
R5238 VDD.n368 VDD.t63 28.5655
R5239 VDD.n368 VDD.t71 28.5655
R5240 VDD.n366 VDD.t59 28.5655
R5241 VDD.n366 VDD.t74 28.5655
R5242 VDD.n364 VDD.t68 28.5655
R5243 VDD.n364 VDD.t65 28.5655
R5244 VDD.n363 VDD.t61 28.5655
R5245 VDD.n363 VDD.t70 28.5655
R5246 VDD.t28 VDD.n123 28.5549
R5247 VDD.n147 VDD.t17 28.5549
R5248 VDD.n299 VDD.t50 27.6484
R5249 VDD.t31 VDD.n267 27.6484
R5250 VDD.t14 VDD.n22 26.7419
R5251 VDD.n154 VDD.t34 26.7419
R5252 VDD.n23 VDD.t20 25.8354
R5253 VDD.t10 VDD.n259 25.8354
R5254 VDD.n304 VDD.n117 25.6005
R5255 VDD.n304 VDD.n303 25.6005
R5256 VDD.n303 VDD.n302 25.6005
R5257 VDD.n302 VDD.n118 25.6005
R5258 VDD.n296 VDD.n118 25.6005
R5259 VDD.n296 VDD.n295 25.6005
R5260 VDD.n295 VDD.n294 25.6005
R5261 VDD.n294 VDD.n125 25.6005
R5262 VDD.n288 VDD.n125 25.6005
R5263 VDD.n288 VDD.n287 25.6005
R5264 VDD.n287 VDD.n286 25.6005
R5265 VDD.n286 VDD.n132 25.6005
R5266 VDD.n280 VDD.n132 25.6005
R5267 VDD.n280 VDD.n279 25.6005
R5268 VDD.n279 VDD.n278 25.6005
R5269 VDD.n278 VDD.n138 25.6005
R5270 VDD.n272 VDD.n138 25.6005
R5271 VDD.n272 VDD.n271 25.6005
R5272 VDD.n271 VDD.n270 25.6005
R5273 VDD.n270 VDD.n145 25.6005
R5274 VDD.n264 VDD.n145 25.6005
R5275 VDD.n264 VDD.n263 25.6005
R5276 VDD.n263 VDD.n262 25.6005
R5277 VDD.n262 VDD.n152 25.6005
R5278 VDD.n255 VDD.n254 25.6005
R5279 VDD.n174 VDD.n171 25.6005
R5280 VDD.n250 VDD.n247 25.6005
R5281 VDD.n247 VDD.n246 25.6005
R5282 VDD.n238 VDD.n235 25.6005
R5283 VDD.n232 VDD.n231 25.6005
R5284 VDD.n228 VDD.n227 25.6005
R5285 VDD.n227 VDD.n224 25.6005
R5286 VDD.n224 VDD.n223 25.6005
R5287 VDD.n223 VDD.n220 25.6005
R5288 VDD.n220 VDD.n219 25.6005
R5289 VDD.n219 VDD.n216 25.6005
R5290 VDD.n215 VDD.n212 25.6005
R5291 VDD.n212 VDD.n211 25.6005
R5292 VDD.n211 VDD.n208 25.6005
R5293 VDD.n208 VDD.n207 25.6005
R5294 VDD.n207 VDD.n205 25.6005
R5295 VDD.n309 VDD.n308 25.6005
R5296 VDD.n308 VDD.n20 25.6005
R5297 VDD.n178 VDD.n20 25.6005
R5298 VDD.n179 VDD.n178 25.6005
R5299 VDD.n180 VDD.n179 25.6005
R5300 VDD.n182 VDD.n180 25.6005
R5301 VDD.n183 VDD.n182 25.6005
R5302 VDD.n184 VDD.n183 25.6005
R5303 VDD.n185 VDD.n184 25.6005
R5304 VDD.n187 VDD.n185 25.6005
R5305 VDD.n188 VDD.n187 25.6005
R5306 VDD.n189 VDD.n188 25.6005
R5307 VDD.n190 VDD.n189 25.6005
R5308 VDD.n192 VDD.n190 25.6005
R5309 VDD.n193 VDD.n192 25.6005
R5310 VDD.n194 VDD.n193 25.6005
R5311 VDD.n195 VDD.n194 25.6005
R5312 VDD.n197 VDD.n195 25.6005
R5313 VDD.n198 VDD.n197 25.6005
R5314 VDD.n199 VDD.n198 25.6005
R5315 VDD.n200 VDD.n199 25.6005
R5316 VDD.n202 VDD.n200 25.6005
R5317 VDD.n203 VDD.n202 25.6005
R5318 VDD.n204 VDD.n203 25.6005
R5319 VDD.n116 VDD.n26 25.6005
R5320 VDD.n27 VDD.n26 25.6005
R5321 VDD.n109 VDD.n27 25.6005
R5322 VDD.n109 VDD.n108 25.6005
R5323 VDD.n108 VDD.n107 25.6005
R5324 VDD.n107 VDD.n29 25.6005
R5325 VDD.n98 VDD.n73 25.6005
R5326 VDD.n93 VDD.n73 25.6005
R5327 VDD.n93 VDD.n92 25.6005
R5328 VDD.n91 VDD.n76 25.6005
R5329 VDD.n86 VDD.n76 25.6005
R5330 VDD.n86 VDD.n85 25.6005
R5331 VDD.n85 VDD.n84 25.6005
R5332 VDD.n84 VDD.n79 25.6005
R5333 VDD.n79 VDD.n12 25.6005
R5334 VDD.n316 VDD.n315 25.6005
R5335 VDD.n315 VDD.n17 25.6005
R5336 VDD.n310 VDD.n17 25.6005
R5337 VDD.n242 VDD.n175 23.3417
R5338 VDD.n102 VDD.n32 21.0829
R5339 VDD.n323 VDD.n322 21.0829
R5340 VDD.n251 VDD.n174 19.577
R5341 VDD.n239 VDD.n238 17.3181
R5342 VDD.n101 VDD.n33 17.3181
R5343 VDD.n318 VDD.n13 17.3181
R5344 VDD.n99 VDD.n98 15.0593
R5345 VDD.n317 VDD.n316 15.0593
R5346 VDD.n235 VDD.n177 14.3064
R5347 VDD.n0 VDD.t21 14.285
R5348 VDD.n254 VDD.n253 13.5534
R5349 VDD.n253 VDD.n171 12.0476
R5350 VDD.n232 VDD.n177 11.2946
R5351 VDD.n99 VDD.n33 10.5417
R5352 VDD.n318 VDD.n317 10.5417
R5353 VDD.n253 VDD.n252 9.43153
R5354 VDD.n240 VDD.n177 9.43153
R5355 VDD.n100 VDD.n99 9.36429
R5356 VDD.n317 VDD.n11 9.36429
R5357 VDD.n252 VDD.n251 9.3005
R5358 VDD.n247 VDD.n172 9.3005
R5359 VDD.n242 VDD.n241 9.3005
R5360 VDD.n240 VDD.n239 9.3005
R5361 VDD.n101 VDD.n100 9.3005
R5362 VDD.n72 VDD.n32 9.3005
R5363 VDD.n13 VDD.n11 9.3005
R5364 VDD.n324 VDD.n323 9.3005
R5365 VDD.n239 VDD.n175 8.28285
R5366 VDD.n32 VDD.n29 8.28285
R5367 VDD.n102 VDD.n101 8.28285
R5368 VDD.n323 VDD.n12 8.28285
R5369 VDD.n322 VDD.n13 8.28285
R5370 VDD.n251 VDD.n250 6.02403
R5371 VDD.n306 VDD.t20 4.98619
R5372 VDD.n260 VDD.t10 4.98619
R5373 VDD.n300 VDD.t14 4.0797
R5374 VDD.n266 VDD.t34 4.0797
R5375 VDD.n72 VDD.n71 3.70853
R5376 VDD.n342 VDD.n324 3.70853
R5377 VDD.t50 VDD.n298 3.17321
R5378 VDD.n268 VDD.t31 3.17321
R5379 VDD.n3 VDD.n1 3.06997
R5380 VDD.n362 VDD.n361 2.73818
R5381 VDD.n342 VDD.n341 2.73818
R5382 VDD.n51 VDD.n50 2.73818
R5383 VDD.n71 VDD.n70 2.73818
R5384 VDD.n373 VDD.n372 2.45598
R5385 VDD.n292 VDD.t28 2.26672
R5386 VDD.n274 VDD.t17 2.26672
R5387 VDD.n243 VDD.n242 2.25932
R5388 VDD.n176 VDD.n10 2.20937
R5389 VDD.n374 VDD.n362 2.07758
R5390 VDD.n376 VDD.n9 1.82938
R5391 VDD.n374 VDD.n373 1.63948
R5392 VDD VDD.n376 1.52224
R5393 VDD.n51 VDD.n10 1.485
R5394 VDD.t5 VDD.n290 1.36023
R5395 VDD.n276 VDD.t2 1.36023
R5396 VDD.n375 VDD.n374 0.9725
R5397 VDD.n5 VDD.n3 0.61449
R5398 VDD.n7 VDD.n5 0.61449
R5399 VDD.n9 VDD.n7 0.61449
R5400 VDD.n71 VDD.n53 0.61449
R5401 VDD.n53 VDD.n51 0.61449
R5402 VDD.n344 VDD.n342 0.61449
R5403 VDD.n362 VDD.n344 0.61449
R5404 VDD.n367 VDD.n365 0.61449
R5405 VDD.n369 VDD.n367 0.61449
R5406 VDD.n373 VDD.n369 0.61449
R5407 VDD.n375 VDD.n10 0.590949
R5408 VDD.n376 VDD.n375 0.4545
R5409 VDD.n284 VDD.t0 0.453744
R5410 VDD.n282 VDD.t7 0.453744
R5411 VDD.n356 VDD.n347 0.38373
R5412 VDD.n351 VDD.n346 0.38373
R5413 VDD.n331 VDD.n330 0.38373
R5414 VDD.n337 VDD.n326 0.38373
R5415 VDD.n45 VDD.n44 0.383729
R5416 VDD.n38 VDD.n35 0.383729
R5417 VDD.n59 VDD.n57 0.383729
R5418 VDD.n66 VDD.n65 0.383729
R5419 VDD.n355 VDD.n348 0.338735
R5420 VDD.n348 VDD.n345 0.338735
R5421 VDD.n361 VDD.n345 0.338735
R5422 VDD.n336 VDD.n327 0.338735
R5423 VDD.n336 VDD.n325 0.338735
R5424 VDD.n341 VDD.n325 0.338735
R5425 VDD.n40 VDD.n36 0.338735
R5426 VDD.n40 VDD.n34 0.338735
R5427 VDD.n50 VDD.n34 0.338735
R5428 VDD.n60 VDD.n55 0.338735
R5429 VDD.n55 VDD.n54 0.338735
R5430 VDD.n70 VDD.n54 0.338735
R5431 VDD.n355 VDD.n354 0.285826
R5432 VDD.n349 VDD.n348 0.285826
R5433 VDD.n328 VDD.n327 0.285826
R5434 VDD.n336 VDD.n335 0.285826
R5435 VDD.n43 VDD.n36 0.285826
R5436 VDD.n41 VDD.n40 0.285826
R5437 VDD.n61 VDD.n60 0.285826
R5438 VDD.n63 VDD.n55 0.285826
R5439 VDD.n351 VDD.n350 0.188
R5440 VDD.n352 VDD.n351 0.188
R5441 VDD.n352 VDD.n347 0.188
R5442 VDD.n353 VDD.n349 0.188
R5443 VDD.n354 VDD.n353 0.188
R5444 VDD.n332 VDD.n331 0.188
R5445 VDD.n332 VDD.n326 0.188
R5446 VDD.n334 VDD.n326 0.188
R5447 VDD.n333 VDD.n328 0.188
R5448 VDD.n335 VDD.n333 0.188
R5449 VDD.n42 VDD.n41 0.188
R5450 VDD.n43 VDD.n42 0.188
R5451 VDD.n39 VDD.n38 0.188
R5452 VDD.n38 VDD.n37 0.188
R5453 VDD.n44 VDD.n37 0.188
R5454 VDD.n62 VDD.n61 0.188
R5455 VDD.n63 VDD.n62 0.188
R5456 VDD.n57 VDD.n56 0.188
R5457 VDD.n65 VDD.n56 0.188
R5458 VDD.n65 VDD.n64 0.188
R5459 VDD.n45 VDD.n36 0.0984044
R5460 VDD.n40 VDD.n35 0.0984044
R5461 VDD.n60 VDD.n59 0.0984044
R5462 VDD.n66 VDD.n55 0.0984044
R5463 VDD.n348 VDD.n346 0.0984028
R5464 VDD.n356 VDD.n355 0.0984028
R5465 VDD.n337 VDD.n336 0.0984028
R5466 VDD.n330 VDD.n327 0.0984028
R5467 VDD.n372 VDD.n371 0.0793043
R5468 VDD.n252 VDD.n172 0.0729138
R5469 VDD.n241 VDD.n240 0.0729138
R5470 VDD.n241 VDD.n176 0.0686034
R5471 VDD.n100 VDD.n72 0.0677414
R5472 VDD.n324 VDD.n11 0.0677414
R5473 VDD.n176 VDD.n172 0.063431
R5474 a_2080_2896.n87 a_2080_2896.n86 185
R5475 a_2080_2896.n86 a_2080_2896.n85 185
R5476 a_2080_2896.n86 a_2080_2896.n8 185
R5477 a_2080_2896.n86 a_2080_2896.n7 185
R5478 a_2080_2896.n86 a_2080_2896.n6 185
R5479 a_2080_2896.n86 a_2080_2896.n5 185
R5480 a_2080_2896.n86 a_2080_2896.n4 185
R5481 a_2080_2896.n53 a_2080_2896.n52 185
R5482 a_2080_2896.n53 a_2080_2896.n40 185
R5483 a_2080_2896.n53 a_2080_2896.n39 185
R5484 a_2080_2896.n53 a_2080_2896.n37 185
R5485 a_2080_2896.n53 a_2080_2896.n36 185
R5486 a_2080_2896.n54 a_2080_2896.n53 185
R5487 a_2080_2896.t2 a_2080_2896.n92 180.167
R5488 a_2080_2896.t2 a_2080_2896.n92 180.167
R5489 a_2080_2896.n21 a_2080_2896.t35 165.607
R5490 a_2080_2896.n9 a_2080_2896.t22 165.607
R5491 a_2080_2896.n70 a_2080_2896.t20 165.032
R5492 a_2080_2896.n19 a_2080_2896.t21 165.032
R5493 a_2080_2896.n18 a_2080_2896.t8 165.032
R5494 a_2080_2896.n17 a_2080_2896.t18 165.032
R5495 a_2080_2896.n16 a_2080_2896.t29 165.032
R5496 a_2080_2896.n15 a_2080_2896.t28 165.032
R5497 a_2080_2896.n14 a_2080_2896.t39 165.032
R5498 a_2080_2896.n13 a_2080_2896.t40 165.032
R5499 a_2080_2896.n12 a_2080_2896.t11 165.032
R5500 a_2080_2896.n11 a_2080_2896.t10 165.032
R5501 a_2080_2896.n10 a_2080_2896.t9 165.032
R5502 a_2080_2896.n9 a_2080_2896.t30 165.032
R5503 a_2080_2896.n68 a_2080_2896.t42 163.058
R5504 a_2080_2896.n66 a_2080_2896.t31 163.058
R5505 a_2080_2896.n64 a_2080_2896.t41 163.058
R5506 a_2080_2896.n62 a_2080_2896.t13 163.058
R5507 a_2080_2896.n60 a_2080_2896.t12 163.058
R5508 a_2080_2896.n32 a_2080_2896.t25 163.058
R5509 a_2080_2896.n58 a_2080_2896.t23 163.058
R5510 a_2080_2896.n28 a_2080_2896.t34 163.058
R5511 a_2080_2896.n26 a_2080_2896.t33 163.058
R5512 a_2080_2896.n24 a_2080_2896.t32 163.058
R5513 a_2080_2896.n22 a_2080_2896.t15 163.058
R5514 a_2080_2896.n20 a_2080_2896.t43 163.058
R5515 a_2080_2896.t3 a_2080_2896.n56 162.941
R5516 a_2080_2896.n56 a_2080_2896.t5 162.941
R5517 a_2080_2896.n68 a_2080_2896.t26 162.781
R5518 a_2080_2896.n66 a_2080_2896.t14 162.781
R5519 a_2080_2896.n64 a_2080_2896.t24 162.781
R5520 a_2080_2896.n62 a_2080_2896.t37 162.781
R5521 a_2080_2896.n60 a_2080_2896.t36 162.781
R5522 a_2080_2896.n28 a_2080_2896.t19 162.781
R5523 a_2080_2896.n26 a_2080_2896.t17 162.781
R5524 a_2080_2896.n24 a_2080_2896.t16 162.781
R5525 a_2080_2896.n22 a_2080_2896.t38 162.781
R5526 a_2080_2896.n20 a_2080_2896.t27 162.781
R5527 a_2080_2896.n57 a_2080_2896.t3 162.639
R5528 a_2080_2896.t5 a_2080_2896.n33 162.639
R5529 a_2080_2896.n91 a_2080_2896.t0 130.75
R5530 a_2080_2896.n86 a_2080_2896.n3 86.5152
R5531 a_2080_2896.n53 a_2080_2896.n38 86.5152
R5532 a_2080_2896.n88 a_2080_2896.n0 30.3012
R5533 a_2080_2896.n73 a_2080_2896.n4 24.8476
R5534 a_2080_2896.n46 a_2080_2896.n39 24.8476
R5535 a_2080_2896.n44 a_2080_2896.n37 24.8476
R5536 a_2080_2896.n75 a_2080_2896.n5 23.3417
R5537 a_2080_2896.n48 a_2080_2896.n40 23.3417
R5538 a_2080_2896.n42 a_2080_2896.n36 23.3417
R5539 a_2080_2896.n72 a_2080_2896.n3 22.0256
R5540 a_2080_2896.n77 a_2080_2896.n6 21.8358
R5541 a_2080_2896.n52 a_2080_2896.n51 21.8358
R5542 a_2080_2896.n54 a_2080_2896.n35 21.8358
R5543 a_2080_2896.n79 a_2080_2896.n7 20.3299
R5544 a_2080_2896.n81 a_2080_2896.n8 18.824
R5545 a_2080_2896.n85 a_2080_2896.n84 17.3181
R5546 a_2080_2896.n86 a_2080_2896.n0 16.3559
R5547 a_2080_2896.n87 a_2080_2896.n2 15.8123
R5548 a_2080_2896.n52 a_2080_2896.n41 14.5711
R5549 a_2080_2896.n55 a_2080_2896.n54 14.5711
R5550 a_2080_2896.n72 a_2080_2896.n71 12.9589
R5551 a_2080_2896.n73 a_2080_2896.n3 12.7256
R5552 a_2080_2896.n46 a_2080_2896.n38 12.7256
R5553 a_2080_2896.n44 a_2080_2896.n38 12.7256
R5554 a_2080_2896.n88 a_2080_2896.n87 11.2946
R5555 a_2080_2896.n85 a_2080_2896.n2 9.78874
R5556 a_2080_2896.n47 a_2080_2896.n46 9.3005
R5557 a_2080_2896.n49 a_2080_2896.n48 9.3005
R5558 a_2080_2896.n51 a_2080_2896.n50 9.3005
R5559 a_2080_2896.n45 a_2080_2896.n44 9.3005
R5560 a_2080_2896.n43 a_2080_2896.n42 9.3005
R5561 a_2080_2896.n35 a_2080_2896.n34 9.3005
R5562 a_2080_2896.n74 a_2080_2896.n73 9.3005
R5563 a_2080_2896.n76 a_2080_2896.n75 9.3005
R5564 a_2080_2896.n78 a_2080_2896.n77 9.3005
R5565 a_2080_2896.n80 a_2080_2896.n79 9.3005
R5566 a_2080_2896.n82 a_2080_2896.n81 9.3005
R5567 a_2080_2896.n84 a_2080_2896.n83 9.3005
R5568 a_2080_2896.n2 a_2080_2896.n1 9.3005
R5569 a_2080_2896.n89 a_2080_2896.n88 9.3005
R5570 a_2080_2896.n71 a_2080_2896.n70 8.61608
R5571 a_2080_2896.n84 a_2080_2896.n8 8.28285
R5572 a_2080_2896.n81 a_2080_2896.n7 6.77697
R5573 a_2080_2896.n53 a_2080_2896.t6 5.8005
R5574 a_2080_2896.n53 a_2080_2896.t4 5.8005
R5575 a_2080_2896.n79 a_2080_2896.n6 5.27109
R5576 a_2080_2896.n77 a_2080_2896.n5 3.76521
R5577 a_2080_2896.n51 a_2080_2896.n40 3.76521
R5578 a_2080_2896.n36 a_2080_2896.n35 3.76521
R5579 a_2080_2896.n86 a_2080_2896.t7 2.48621
R5580 a_2080_2896.n86 a_2080_2896.t1 2.48621
R5581 a_2080_2896.n90 a_2080_2896.n0 2.36936
R5582 a_2080_2896.n75 a_2080_2896.n4 2.25932
R5583 a_2080_2896.n48 a_2080_2896.n39 2.25932
R5584 a_2080_2896.n42 a_2080_2896.n37 2.25932
R5585 a_2080_2896.n69 a_2080_2896.n68 2.25162
R5586 a_2080_2896.n67 a_2080_2896.n66 2.25162
R5587 a_2080_2896.n65 a_2080_2896.n64 2.25162
R5588 a_2080_2896.n63 a_2080_2896.n62 2.25162
R5589 a_2080_2896.n61 a_2080_2896.n60 2.25162
R5590 a_2080_2896.n32 a_2080_2896.n30 2.25162
R5591 a_2080_2896.n59 a_2080_2896.n58 2.25162
R5592 a_2080_2896.n29 a_2080_2896.n28 2.25162
R5593 a_2080_2896.n27 a_2080_2896.n26 2.25162
R5594 a_2080_2896.n25 a_2080_2896.n24 2.25162
R5595 a_2080_2896.n23 a_2080_2896.n22 2.25162
R5596 a_2080_2896.n21 a_2080_2896.n20 2.25162
R5597 a_2080_2896.n71 a_2080_2896.n19 2.17137
R5598 a_2080_2896.n92 a_2080_2896.n91 1.27148
R5599 a_2080_2896.n23 a_2080_2896.n21 0.574917
R5600 a_2080_2896.n25 a_2080_2896.n23 0.574917
R5601 a_2080_2896.n27 a_2080_2896.n25 0.574917
R5602 a_2080_2896.n29 a_2080_2896.n27 0.574917
R5603 a_2080_2896.n30 a_2080_2896.n29 0.574917
R5604 a_2080_2896.n59 a_2080_2896.n30 0.574917
R5605 a_2080_2896.n61 a_2080_2896.n59 0.574917
R5606 a_2080_2896.n63 a_2080_2896.n61 0.574917
R5607 a_2080_2896.n65 a_2080_2896.n63 0.574917
R5608 a_2080_2896.n67 a_2080_2896.n65 0.574917
R5609 a_2080_2896.n69 a_2080_2896.n67 0.574917
R5610 a_2080_2896.n70 a_2080_2896.n69 0.574917
R5611 a_2080_2896.n10 a_2080_2896.n9 0.574917
R5612 a_2080_2896.n11 a_2080_2896.n10 0.574917
R5613 a_2080_2896.n12 a_2080_2896.n11 0.574917
R5614 a_2080_2896.n13 a_2080_2896.n12 0.574917
R5615 a_2080_2896.n14 a_2080_2896.n13 0.574917
R5616 a_2080_2896.n15 a_2080_2896.n14 0.574917
R5617 a_2080_2896.n16 a_2080_2896.n15 0.574917
R5618 a_2080_2896.n17 a_2080_2896.n16 0.574917
R5619 a_2080_2896.n18 a_2080_2896.n17 0.574917
R5620 a_2080_2896.n19 a_2080_2896.n18 0.574917
R5621 a_2080_2896.n91 a_2080_2896.n90 0.320353
R5622 a_2080_2896.n33 a_2080_2896.n31 0.302413
R5623 a_2080_2896.n57 a_2080_2896.n31 0.302413
R5624 a_2080_2896.n41 a_2080_2896.n31 0.217891
R5625 a_2080_2896.n56 a_2080_2896.n55 0.217891
R5626 a_2080_2896.n50 a_2080_2896.n41 0.196152
R5627 a_2080_2896.n50 a_2080_2896.n49 0.196152
R5628 a_2080_2896.n49 a_2080_2896.n47 0.196152
R5629 a_2080_2896.n47 a_2080_2896.n45 0.196152
R5630 a_2080_2896.n45 a_2080_2896.n43 0.196152
R5631 a_2080_2896.n43 a_2080_2896.n34 0.196152
R5632 a_2080_2896.n55 a_2080_2896.n34 0.196152
R5633 a_2080_2896.n90 a_2080_2896.n89 0.196152
R5634 a_2080_2896.n89 a_2080_2896.n1 0.196152
R5635 a_2080_2896.n83 a_2080_2896.n1 0.196152
R5636 a_2080_2896.n83 a_2080_2896.n82 0.196152
R5637 a_2080_2896.n82 a_2080_2896.n80 0.196152
R5638 a_2080_2896.n80 a_2080_2896.n78 0.196152
R5639 a_2080_2896.n78 a_2080_2896.n76 0.196152
R5640 a_2080_2896.n76 a_2080_2896.n74 0.196152
R5641 a_2080_2896.n74 a_2080_2896.n72 0.196152
R5642 a_2080_2896.n33 a_2080_2896.n32 0.142018
R5643 a_2080_2896.n58 a_2080_2896.n57 0.142018
R5644 a_4920_2896.n46 a_4920_2896.n28 185
R5645 a_4920_2896.n46 a_4920_2896.n27 185
R5646 a_4920_2896.n46 a_4920_2896.n26 185
R5647 a_4920_2896.n46 a_4920_2896.n25 185
R5648 a_4920_2896.n46 a_4920_2896.n24 185
R5649 a_4920_2896.n46 a_4920_2896.n23 185
R5650 a_4920_2896.n46 a_4920_2896.n22 185
R5651 a_4920_2896.n30 a_4920_2896.t25 130.75
R5652 a_4920_2896.n30 a_4920_2896.t26 91.3557
R5653 a_4920_2896.n47 a_4920_2896.n46 86.5152
R5654 a_4920_2896.n45 a_4920_2896.n29 30.3012
R5655 a_4920_2896.n15 a_4920_2896.n14 26.8581
R5656 a_4920_2896.n5 a_4920_2896.n4 26.6299
R5657 a_4920_2896.n19 a_4920_2896.n9 25.7063
R5658 a_4920_2896.n18 a_4920_2896.n10 25.7063
R5659 a_4920_2896.n17 a_4920_2896.n11 25.7063
R5660 a_4920_2896.n16 a_4920_2896.n12 25.7063
R5661 a_4920_2896.n15 a_4920_2896.n13 25.7063
R5662 a_4920_2896.n51 a_4920_2896.n50 25.4783
R5663 a_4920_2896.n5 a_4920_2896.n3 25.4781
R5664 a_4920_2896.n6 a_4920_2896.n2 25.4781
R5665 a_4920_2896.n7 a_4920_2896.n1 25.4781
R5666 a_4920_2896.n8 a_4920_2896.n0 25.4781
R5667 a_4920_2896.n22 a_4920_2896.n21 24.8476
R5668 a_4920_2896.n31 a_4920_2896.n23 23.3417
R5669 a_4920_2896.n48 a_4920_2896.n47 22.0256
R5670 a_4920_2896.n33 a_4920_2896.n24 21.8358
R5671 a_4920_2896.n35 a_4920_2896.n25 20.3299
R5672 a_4920_2896.n37 a_4920_2896.n26 18.824
R5673 a_4920_2896.n39 a_4920_2896.n27 17.3181
R5674 a_4920_2896.n46 a_4920_2896.n45 16.3559
R5675 a_4920_2896.n41 a_4920_2896.n28 15.8123
R5676 a_4920_2896.n47 a_4920_2896.n21 12.7256
R5677 a_4920_2896.n29 a_4920_2896.n28 11.2946
R5678 a_4920_2896.n41 a_4920_2896.n27 9.78874
R5679 a_4920_2896.n49 a_4920_2896.n19 9.30285
R5680 a_4920_2896.n21 a_4920_2896.n20 9.3005
R5681 a_4920_2896.n32 a_4920_2896.n31 9.3005
R5682 a_4920_2896.n34 a_4920_2896.n33 9.3005
R5683 a_4920_2896.n36 a_4920_2896.n35 9.3005
R5684 a_4920_2896.n38 a_4920_2896.n37 9.3005
R5685 a_4920_2896.n40 a_4920_2896.n39 9.3005
R5686 a_4920_2896.n42 a_4920_2896.n41 9.3005
R5687 a_4920_2896.n43 a_4920_2896.n29 9.3005
R5688 a_4920_2896.n39 a_4920_2896.n26 8.28285
R5689 a_4920_2896.n37 a_4920_2896.n25 6.77697
R5690 a_4920_2896.n4 a_4920_2896.t14 5.8005
R5691 a_4920_2896.n4 a_4920_2896.t9 5.8005
R5692 a_4920_2896.n3 a_4920_2896.t22 5.8005
R5693 a_4920_2896.n3 a_4920_2896.t21 5.8005
R5694 a_4920_2896.n2 a_4920_2896.t20 5.8005
R5695 a_4920_2896.n2 a_4920_2896.t3 5.8005
R5696 a_4920_2896.n1 a_4920_2896.t4 5.8005
R5697 a_4920_2896.n1 a_4920_2896.t11 5.8005
R5698 a_4920_2896.n0 a_4920_2896.t10 5.8005
R5699 a_4920_2896.n0 a_4920_2896.t16 5.8005
R5700 a_4920_2896.n9 a_4920_2896.t8 5.8005
R5701 a_4920_2896.n9 a_4920_2896.t1 5.8005
R5702 a_4920_2896.n10 a_4920_2896.t18 5.8005
R5703 a_4920_2896.n10 a_4920_2896.t2 5.8005
R5704 a_4920_2896.n11 a_4920_2896.t13 5.8005
R5705 a_4920_2896.n11 a_4920_2896.t19 5.8005
R5706 a_4920_2896.n12 a_4920_2896.t5 5.8005
R5707 a_4920_2896.n12 a_4920_2896.t12 5.8005
R5708 a_4920_2896.n13 a_4920_2896.t7 5.8005
R5709 a_4920_2896.n13 a_4920_2896.t6 5.8005
R5710 a_4920_2896.n14 a_4920_2896.t0 5.8005
R5711 a_4920_2896.n14 a_4920_2896.t17 5.8005
R5712 a_4920_2896.t23 a_4920_2896.n51 5.8005
R5713 a_4920_2896.n51 a_4920_2896.t15 5.8005
R5714 a_4920_2896.n35 a_4920_2896.n24 5.27109
R5715 a_4920_2896.n33 a_4920_2896.n23 3.76521
R5716 a_4920_2896.n50 a_4920_2896.n49 2.92217
R5717 a_4920_2896.n46 a_4920_2896.t26 2.48621
R5718 a_4920_2896.n46 a_4920_2896.t24 2.48621
R5719 a_4920_2896.n45 a_4920_2896.n44 2.36936
R5720 a_4920_2896.n31 a_4920_2896.n22 2.25932
R5721 a_4920_2896.n49 a_4920_2896.n48 2.19829
R5722 a_4920_2896.n16 a_4920_2896.n15 1.15229
R5723 a_4920_2896.n17 a_4920_2896.n16 1.15229
R5724 a_4920_2896.n18 a_4920_2896.n17 1.15229
R5725 a_4920_2896.n19 a_4920_2896.n18 1.15229
R5726 a_4920_2896.n6 a_4920_2896.n5 1.15229
R5727 a_4920_2896.n7 a_4920_2896.n6 1.15229
R5728 a_4920_2896.n8 a_4920_2896.n7 1.15229
R5729 a_4920_2896.n50 a_4920_2896.n8 1.15229
R5730 a_4920_2896.n44 a_4920_2896.n30 0.320353
R5731 a_4920_2896.n44 a_4920_2896.n43 0.196152
R5732 a_4920_2896.n43 a_4920_2896.n42 0.196152
R5733 a_4920_2896.n42 a_4920_2896.n40 0.196152
R5734 a_4920_2896.n40 a_4920_2896.n38 0.196152
R5735 a_4920_2896.n38 a_4920_2896.n36 0.196152
R5736 a_4920_2896.n36 a_4920_2896.n34 0.196152
R5737 a_4920_2896.n34 a_4920_2896.n32 0.196152
R5738 a_4920_2896.n32 a_4920_2896.n20 0.196152
R5739 a_4920_2896.n48 a_4920_2896.n20 0.196152
R5740 VP.n0 VP.t7 263.647
R5741 VP.n3 VP.t3 262.863
R5742 VP.n2 VP.t1 262.498
R5743 VP.n0 VP.t6 261.709
R5744 VP.n1 VP.t2 261.709
R5745 VP.n3 VP.t5 261.584
R5746 VP.n4 VP.t4 261.584
R5747 VP.n5 VP.t0 261.433
R5748 VP.n6 VP.n2 8.91083
R5749 VP VP.n6 2.38312
R5750 VP.n1 VP.n0 1.72698
R5751 VP.n6 VP.n5 1.52193
R5752 VP.n5 VP.n4 1.4312
R5753 VP.n4 VP.n3 1.16675
R5754 VP.n2 VP.n1 1.14999
R5755 a_2995_7336.n32 a_2995_7336.n31 185
R5756 a_2995_7336.n32 a_2995_7336.n14 185
R5757 a_2995_7336.n32 a_2995_7336.n13 185
R5758 a_2995_7336.n32 a_2995_7336.n12 185
R5759 a_2995_7336.n32 a_2995_7336.n11 185
R5760 a_2995_7336.n32 a_2995_7336.n10 185
R5761 a_2995_7336.n32 a_2995_7336.n9 185
R5762 a_2995_7336.n15 a_2995_7336.t17 130.75
R5763 a_2995_7336.n15 a_2995_7336.t19 91.3557
R5764 a_2995_7336.n33 a_2995_7336.n32 86.5152
R5765 a_2995_7336.n17 a_2995_7336.n8 30.3012
R5766 a_2995_7336.n31 a_2995_7336.n7 24.8476
R5767 a_2995_7336.n30 a_2995_7336.n14 23.3417
R5768 a_2995_7336.n34 a_2995_7336.n33 22.0256
R5769 a_2995_7336.n27 a_2995_7336.n13 21.8358
R5770 a_2995_7336.n25 a_2995_7336.n12 20.3299
R5771 a_2995_7336.n23 a_2995_7336.n11 18.824
R5772 a_2995_7336.n21 a_2995_7336.n10 17.3181
R5773 a_2995_7336.n32 a_2995_7336.n8 16.3559
R5774 a_2995_7336.n19 a_2995_7336.n9 15.8123
R5775 a_2995_7336.n33 a_2995_7336.n7 12.7256
R5776 a_2995_7336.n38 a_2995_7336.n37 12.1709
R5777 a_2995_7336.n39 a_2995_7336.n38 12.1709
R5778 a_2995_7336.n40 a_2995_7336.n0 11.493
R5779 a_2995_7336.n37 a_2995_7336.n35 11.493
R5780 a_2995_7336.n3 a_2995_7336.n1 11.493
R5781 a_2995_7336.n39 a_2995_7336.n4 11.493
R5782 a_2995_7336.n41 a_2995_7336.n40 11.493
R5783 a_2995_7336.n37 a_2995_7336.n36 11.4929
R5784 a_2995_7336.n3 a_2995_7336.n2 11.4929
R5785 a_2995_7336.n39 a_2995_7336.n5 11.4929
R5786 a_2995_7336.n17 a_2995_7336.n9 11.2946
R5787 a_2995_7336.n19 a_2995_7336.n10 9.78874
R5788 a_2995_7336.n7 a_2995_7336.n6 9.3005
R5789 a_2995_7336.n30 a_2995_7336.n29 9.3005
R5790 a_2995_7336.n28 a_2995_7336.n27 9.3005
R5791 a_2995_7336.n26 a_2995_7336.n25 9.3005
R5792 a_2995_7336.n24 a_2995_7336.n23 9.3005
R5793 a_2995_7336.n22 a_2995_7336.n21 9.3005
R5794 a_2995_7336.n20 a_2995_7336.n19 9.3005
R5795 a_2995_7336.n18 a_2995_7336.n17 9.3005
R5796 a_2995_7336.n21 a_2995_7336.n11 8.28285
R5797 a_2995_7336.n23 a_2995_7336.n12 6.77697
R5798 a_2995_7336.n25 a_2995_7336.n13 5.27109
R5799 a_2995_7336.n27 a_2995_7336.n14 3.76521
R5800 a_2995_7336.n38 a_2995_7336.n34 3.48602
R5801 a_2995_7336.n0 a_2995_7336.t3 2.48621
R5802 a_2995_7336.n0 a_2995_7336.t8 2.48621
R5803 a_2995_7336.n36 a_2995_7336.t14 2.48621
R5804 a_2995_7336.n36 a_2995_7336.t2 2.48621
R5805 a_2995_7336.n35 a_2995_7336.t16 2.48621
R5806 a_2995_7336.n35 a_2995_7336.t13 2.48621
R5807 a_2995_7336.n2 a_2995_7336.t6 2.48621
R5808 a_2995_7336.n2 a_2995_7336.t10 2.48621
R5809 a_2995_7336.n1 a_2995_7336.t12 2.48621
R5810 a_2995_7336.n1 a_2995_7336.t5 2.48621
R5811 a_2995_7336.n5 a_2995_7336.t4 2.48621
R5812 a_2995_7336.n5 a_2995_7336.t11 2.48621
R5813 a_2995_7336.n4 a_2995_7336.t7 2.48621
R5814 a_2995_7336.n4 a_2995_7336.t15 2.48621
R5815 a_2995_7336.n32 a_2995_7336.t1 2.48621
R5816 a_2995_7336.n32 a_2995_7336.t18 2.48621
R5817 a_2995_7336.n41 a_2995_7336.t9 2.48621
R5818 a_2995_7336.t0 a_2995_7336.n41 2.48621
R5819 a_2995_7336.n16 a_2995_7336.n8 2.36936
R5820 a_2995_7336.n31 a_2995_7336.n30 2.25932
R5821 a_2995_7336.n37 a_2995_7336.n3 1.15229
R5822 a_2995_7336.n40 a_2995_7336.n3 1.15229
R5823 a_2995_7336.n40 a_2995_7336.n39 1.15229
R5824 a_2995_7336.n16 a_2995_7336.n15 0.320353
R5825 a_2995_7336.n34 a_2995_7336.n6 0.196152
R5826 a_2995_7336.n29 a_2995_7336.n6 0.196152
R5827 a_2995_7336.n29 a_2995_7336.n28 0.196152
R5828 a_2995_7336.n28 a_2995_7336.n26 0.196152
R5829 a_2995_7336.n26 a_2995_7336.n24 0.196152
R5830 a_2995_7336.n24 a_2995_7336.n22 0.196152
R5831 a_2995_7336.n22 a_2995_7336.n20 0.196152
R5832 a_2995_7336.n20 a_2995_7336.n18 0.196152
R5833 a_2995_7336.n18 a_2995_7336.n16 0.196152
R5834 VN.n0 VN.t0 263.647
R5835 VN.n3 VN.t2 262.863
R5836 VN.n2 VN.t5 262.498
R5837 VN.n1 VN.t4 261.709
R5838 VN.n0 VN.t1 261.709
R5839 VN.n4 VN.t7 261.584
R5840 VN.n3 VN.t6 261.584
R5841 VN.n5 VN.t3 261.433
R5842 VN.n6 VN.n2 8.91083
R5843 VN VN.n6 2.48729
R5844 VN.n1 VN.n0 1.72698
R5845 VN.n6 VN.n5 1.52193
R5846 VN.n5 VN.n4 1.4312
R5847 VN.n4 VN.n3 1.16675
R5848 VN.n2 VN.n1 1.14999
R5849 a_2479_9004.n70 a_2479_9004.t22 260.111
R5850 a_2479_9004.n4 a_2479_9004.t21 260.111
R5851 a_2479_9004.n3 a_2479_9004.t0 260.111
R5852 a_2479_9004.n1 a_2479_9004.t2 260.111
R5853 a_2479_9004.n70 a_2479_9004.t4 260.111
R5854 a_2479_9004.n4 a_2479_9004.t6 260.111
R5855 a_2479_9004.n3 a_2479_9004.t24 260.111
R5856 a_2479_9004.n1 a_2479_9004.t23 260.111
R5857 a_2479_9004.n2 a_2479_9004.n0 203.413
R5858 a_2479_9004.n72 a_2479_9004.n71 203.412
R5859 a_2479_9004.n34 a_2479_9004.n33 185
R5860 a_2479_9004.n34 a_2479_9004.n16 185
R5861 a_2479_9004.n34 a_2479_9004.n15 185
R5862 a_2479_9004.n34 a_2479_9004.n14 185
R5863 a_2479_9004.n34 a_2479_9004.n13 185
R5864 a_2479_9004.n34 a_2479_9004.n12 185
R5865 a_2479_9004.n34 a_2479_9004.n11 185
R5866 a_2479_9004.n65 a_2479_9004.n64 185
R5867 a_2479_9004.n65 a_2479_9004.n47 185
R5868 a_2479_9004.n65 a_2479_9004.n46 185
R5869 a_2479_9004.n65 a_2479_9004.n45 185
R5870 a_2479_9004.n65 a_2479_9004.n44 185
R5871 a_2479_9004.n65 a_2479_9004.n43 185
R5872 a_2479_9004.n65 a_2479_9004.n42 185
R5873 a_2479_9004.n17 a_2479_9004.t8 130.75
R5874 a_2479_9004.n48 a_2479_9004.t11 130.75
R5875 a_2479_9004.n17 a_2479_9004.t10 91.3557
R5876 a_2479_9004.n48 a_2479_9004.t12 91.3557
R5877 a_2479_9004.n35 a_2479_9004.n34 86.5152
R5878 a_2479_9004.n66 a_2479_9004.n65 86.5152
R5879 a_2479_9004.n19 a_2479_9004.n10 30.3012
R5880 a_2479_9004.n50 a_2479_9004.n41 30.3012
R5881 a_2479_9004.n0 a_2479_9004.t3 28.5655
R5882 a_2479_9004.n0 a_2479_9004.t1 28.5655
R5883 a_2479_9004.t7 a_2479_9004.n72 28.5655
R5884 a_2479_9004.n72 a_2479_9004.t5 28.5655
R5885 a_2479_9004.n33 a_2479_9004.n9 24.8476
R5886 a_2479_9004.n64 a_2479_9004.n40 24.8476
R5887 a_2479_9004.n32 a_2479_9004.n16 23.3417
R5888 a_2479_9004.n63 a_2479_9004.n47 23.3417
R5889 a_2479_9004.n36 a_2479_9004.n35 22.0256
R5890 a_2479_9004.n67 a_2479_9004.n66 22.0256
R5891 a_2479_9004.n29 a_2479_9004.n15 21.8358
R5892 a_2479_9004.n60 a_2479_9004.n46 21.8358
R5893 a_2479_9004.n27 a_2479_9004.n14 20.3299
R5894 a_2479_9004.n58 a_2479_9004.n45 20.3299
R5895 a_2479_9004.n25 a_2479_9004.n13 18.824
R5896 a_2479_9004.n56 a_2479_9004.n44 18.824
R5897 a_2479_9004.n7 a_2479_9004.n5 17.4823
R5898 a_2479_9004.n23 a_2479_9004.n12 17.3181
R5899 a_2479_9004.n54 a_2479_9004.n43 17.3181
R5900 a_2479_9004.n34 a_2479_9004.n10 16.3559
R5901 a_2479_9004.n65 a_2479_9004.n41 16.3559
R5902 a_2479_9004.n21 a_2479_9004.n11 15.8123
R5903 a_2479_9004.n52 a_2479_9004.n42 15.8123
R5904 a_2479_9004.n7 a_2479_9004.n6 14.6053
R5905 a_2479_9004.n38 a_2479_9004.n37 14.377
R5906 a_2479_9004.n35 a_2479_9004.n9 12.7256
R5907 a_2479_9004.n66 a_2479_9004.n40 12.7256
R5908 a_2479_9004.n19 a_2479_9004.n11 11.2946
R5909 a_2479_9004.n50 a_2479_9004.n42 11.2946
R5910 a_2479_9004.n69 a_2479_9004.n7 10.4849
R5911 a_2479_9004.n21 a_2479_9004.n12 9.78874
R5912 a_2479_9004.n52 a_2479_9004.n43 9.78874
R5913 a_2479_9004.n9 a_2479_9004.n8 9.3005
R5914 a_2479_9004.n32 a_2479_9004.n31 9.3005
R5915 a_2479_9004.n30 a_2479_9004.n29 9.3005
R5916 a_2479_9004.n28 a_2479_9004.n27 9.3005
R5917 a_2479_9004.n26 a_2479_9004.n25 9.3005
R5918 a_2479_9004.n24 a_2479_9004.n23 9.3005
R5919 a_2479_9004.n22 a_2479_9004.n21 9.3005
R5920 a_2479_9004.n20 a_2479_9004.n19 9.3005
R5921 a_2479_9004.n40 a_2479_9004.n39 9.3005
R5922 a_2479_9004.n63 a_2479_9004.n62 9.3005
R5923 a_2479_9004.n61 a_2479_9004.n60 9.3005
R5924 a_2479_9004.n59 a_2479_9004.n58 9.3005
R5925 a_2479_9004.n57 a_2479_9004.n56 9.3005
R5926 a_2479_9004.n55 a_2479_9004.n54 9.3005
R5927 a_2479_9004.n53 a_2479_9004.n52 9.3005
R5928 a_2479_9004.n51 a_2479_9004.n50 9.3005
R5929 a_2479_9004.n70 a_2479_9004.n69 8.69704
R5930 a_2479_9004.n23 a_2479_9004.n13 8.28285
R5931 a_2479_9004.n54 a_2479_9004.n44 8.28285
R5932 a_2479_9004.n25 a_2479_9004.n14 6.77697
R5933 a_2479_9004.n56 a_2479_9004.n45 6.77697
R5934 a_2479_9004.n38 a_2479_9004.n36 6.19091
R5935 a_2479_9004.n27 a_2479_9004.n15 5.27109
R5936 a_2479_9004.n58 a_2479_9004.n46 5.27109
R5937 a_2479_9004.n29 a_2479_9004.n16 3.76521
R5938 a_2479_9004.n60 a_2479_9004.n47 3.76521
R5939 a_2479_9004.n68 a_2479_9004.n67 3.31388
R5940 a_2479_9004.n5 a_2479_9004.t16 2.48621
R5941 a_2479_9004.n5 a_2479_9004.t15 2.48621
R5942 a_2479_9004.n6 a_2479_9004.t20 2.48621
R5943 a_2479_9004.n6 a_2479_9004.t19 2.48621
R5944 a_2479_9004.n34 a_2479_9004.t17 2.48621
R5945 a_2479_9004.n34 a_2479_9004.t9 2.48621
R5946 a_2479_9004.n37 a_2479_9004.t14 2.48621
R5947 a_2479_9004.n37 a_2479_9004.t13 2.48621
R5948 a_2479_9004.n65 a_2479_9004.t12 2.48621
R5949 a_2479_9004.n65 a_2479_9004.t18 2.48621
R5950 a_2479_9004.n18 a_2479_9004.n10 2.36936
R5951 a_2479_9004.n49 a_2479_9004.n41 2.36936
R5952 a_2479_9004.n68 a_2479_9004.n38 2.30287
R5953 a_2479_9004.n33 a_2479_9004.n32 2.25932
R5954 a_2479_9004.n64 a_2479_9004.n63 2.25932
R5955 a_2479_9004.n69 a_2479_9004.n68 1.07418
R5956 a_2479_9004.n18 a_2479_9004.n17 0.320353
R5957 a_2479_9004.n49 a_2479_9004.n48 0.320353
R5958 a_2479_9004.n36 a_2479_9004.n8 0.196152
R5959 a_2479_9004.n31 a_2479_9004.n8 0.196152
R5960 a_2479_9004.n31 a_2479_9004.n30 0.196152
R5961 a_2479_9004.n30 a_2479_9004.n28 0.196152
R5962 a_2479_9004.n28 a_2479_9004.n26 0.196152
R5963 a_2479_9004.n26 a_2479_9004.n24 0.196152
R5964 a_2479_9004.n24 a_2479_9004.n22 0.196152
R5965 a_2479_9004.n22 a_2479_9004.n20 0.196152
R5966 a_2479_9004.n20 a_2479_9004.n18 0.196152
R5967 a_2479_9004.n67 a_2479_9004.n39 0.196152
R5968 a_2479_9004.n62 a_2479_9004.n39 0.196152
R5969 a_2479_9004.n62 a_2479_9004.n61 0.196152
R5970 a_2479_9004.n61 a_2479_9004.n59 0.196152
R5971 a_2479_9004.n59 a_2479_9004.n57 0.196152
R5972 a_2479_9004.n57 a_2479_9004.n55 0.196152
R5973 a_2479_9004.n55 a_2479_9004.n53 0.196152
R5974 a_2479_9004.n53 a_2479_9004.n51 0.196152
R5975 a_2479_9004.n51 a_2479_9004.n49 0.196152
R5976 a_2479_9004.n4 a_2479_9004.n3 0.0850588
R5977 a_2479_9004.n2 a_2479_9004.n1 0.0427794
R5978 a_2479_9004.n3 a_2479_9004.n2 0.0427794
R5979 a_2479_9004.n71 a_2479_9004.n4 0.0427794
R5980 a_2479_9004.n71 a_2479_9004.n70 0.0427794
R5981 a_3758_2896.n33 a_3758_2896.n32 185
R5982 a_3758_2896.n33 a_3758_2896.n15 185
R5983 a_3758_2896.n33 a_3758_2896.n14 185
R5984 a_3758_2896.n33 a_3758_2896.n13 185
R5985 a_3758_2896.n33 a_3758_2896.n12 185
R5986 a_3758_2896.n33 a_3758_2896.n11 185
R5987 a_3758_2896.n33 a_3758_2896.n10 185
R5988 a_3758_2896.n16 a_3758_2896.t13 130.75
R5989 a_3758_2896.n16 a_3758_2896.t14 91.3557
R5990 a_3758_2896.n34 a_3758_2896.n33 86.5152
R5991 a_3758_2896.n18 a_3758_2896.n9 30.3012
R5992 a_3758_2896.n2 a_3758_2896.n0 29.1073
R5993 a_3758_2896.n39 a_3758_2896.n38 27.9576
R5994 a_3758_2896.n37 a_3758_2896.n36 27.9576
R5995 a_3758_2896.n6 a_3758_2896.n5 27.9576
R5996 a_3758_2896.n4 a_3758_2896.n3 27.9576
R5997 a_3758_2896.n2 a_3758_2896.n1 27.9576
R5998 a_3758_2896.n32 a_3758_2896.n8 24.8476
R5999 a_3758_2896.n31 a_3758_2896.n15 23.3417
R6000 a_3758_2896.n35 a_3758_2896.n34 22.0256
R6001 a_3758_2896.n28 a_3758_2896.n14 21.8358
R6002 a_3758_2896.n26 a_3758_2896.n13 20.3299
R6003 a_3758_2896.n24 a_3758_2896.n12 18.824
R6004 a_3758_2896.n22 a_3758_2896.n11 17.3181
R6005 a_3758_2896.n33 a_3758_2896.n9 16.3559
R6006 a_3758_2896.n20 a_3758_2896.n10 15.8123
R6007 a_3758_2896.n34 a_3758_2896.n8 12.7256
R6008 a_3758_2896.n37 a_3758_2896.n35 12.0517
R6009 a_3758_2896.n18 a_3758_2896.n10 11.2946
R6010 a_3758_2896.n20 a_3758_2896.n11 9.78874
R6011 a_3758_2896.n8 a_3758_2896.n7 9.3005
R6012 a_3758_2896.n31 a_3758_2896.n30 9.3005
R6013 a_3758_2896.n29 a_3758_2896.n28 9.3005
R6014 a_3758_2896.n27 a_3758_2896.n26 9.3005
R6015 a_3758_2896.n25 a_3758_2896.n24 9.3005
R6016 a_3758_2896.n23 a_3758_2896.n22 9.3005
R6017 a_3758_2896.n21 a_3758_2896.n20 9.3005
R6018 a_3758_2896.n19 a_3758_2896.n18 9.3005
R6019 a_3758_2896.n22 a_3758_2896.n12 8.28285
R6020 a_3758_2896.n24 a_3758_2896.n13 6.77697
R6021 a_3758_2896.n36 a_3758_2896.t5 5.8005
R6022 a_3758_2896.n36 a_3758_2896.t7 5.8005
R6023 a_3758_2896.n5 a_3758_2896.t2 5.8005
R6024 a_3758_2896.n5 a_3758_2896.t1 5.8005
R6025 a_3758_2896.n3 a_3758_2896.t9 5.8005
R6026 a_3758_2896.n3 a_3758_2896.t8 5.8005
R6027 a_3758_2896.n1 a_3758_2896.t0 5.8005
R6028 a_3758_2896.n1 a_3758_2896.t10 5.8005
R6029 a_3758_2896.n0 a_3758_2896.t3 5.8005
R6030 a_3758_2896.n0 a_3758_2896.t4 5.8005
R6031 a_3758_2896.n39 a_3758_2896.t6 5.8005
R6032 a_3758_2896.t11 a_3758_2896.n39 5.8005
R6033 a_3758_2896.n26 a_3758_2896.n14 5.27109
R6034 a_3758_2896.n28 a_3758_2896.n15 3.76521
R6035 a_3758_2896.n33 a_3758_2896.t14 2.48621
R6036 a_3758_2896.n33 a_3758_2896.t12 2.48621
R6037 a_3758_2896.n17 a_3758_2896.n9 2.36936
R6038 a_3758_2896.n6 a_3758_2896.n4 2.30199
R6039 a_3758_2896.n32 a_3758_2896.n31 2.25932
R6040 a_3758_2896.n4 a_3758_2896.n2 1.1502
R6041 a_3758_2896.n38 a_3758_2896.n6 1.1502
R6042 a_3758_2896.n38 a_3758_2896.n37 1.1502
R6043 a_3758_2896.n17 a_3758_2896.n16 0.320353
R6044 a_3758_2896.n35 a_3758_2896.n7 0.196152
R6045 a_3758_2896.n30 a_3758_2896.n7 0.196152
R6046 a_3758_2896.n30 a_3758_2896.n29 0.196152
R6047 a_3758_2896.n29 a_3758_2896.n27 0.196152
R6048 a_3758_2896.n27 a_3758_2896.n25 0.196152
R6049 a_3758_2896.n25 a_3758_2896.n23 0.196152
R6050 a_3758_2896.n23 a_3758_2896.n21 0.196152
R6051 a_3758_2896.n21 a_3758_2896.n19 0.196152
R6052 a_3758_2896.n19 a_3758_2896.n17 0.196152
R6053 EN.n0 EN.t0 262.997
R6054 EN.n1 EN.t1 262.007
R6055 EN.n0 EN.t2 262.007
R6056 EN.n1 EN.n0 0.989232
R6057 EN EN.n1 0.365614
R6058 C1 C1.t0 17.7454
R6059 C1 C1.t1 0.00167066
R6060 IBIAS.n26 IBIAS.n25 185
R6061 IBIAS.n26 IBIAS.n8 185
R6062 IBIAS.n26 IBIAS.n7 185
R6063 IBIAS.n26 IBIAS.n6 185
R6064 IBIAS.n26 IBIAS.n5 185
R6065 IBIAS.n26 IBIAS.n4 185
R6066 IBIAS.n26 IBIAS.n3 185
R6067 IBIAS.n9 IBIAS.t0 130.75
R6068 IBIAS.n9 IBIAS.t1 91.3557
R6069 IBIAS.n27 IBIAS.n26 86.5152
R6070 IBIAS.n11 IBIAS.n2 30.3012
R6071 IBIAS.n25 IBIAS.n1 24.8476
R6072 IBIAS.n24 IBIAS.n8 23.3417
R6073 IBIAS.n28 IBIAS.n27 22.0256
R6074 IBIAS.n21 IBIAS.n7 21.8358
R6075 IBIAS.n19 IBIAS.n6 20.3299
R6076 IBIAS.n17 IBIAS.n5 18.824
R6077 IBIAS.n15 IBIAS.n4 17.3181
R6078 IBIAS.n26 IBIAS.n2 16.3559
R6079 IBIAS.n13 IBIAS.n3 15.8123
R6080 IBIAS.n27 IBIAS.n1 12.7256
R6081 IBIAS.n11 IBIAS.n3 11.2946
R6082 IBIAS.n13 IBIAS.n4 9.78874
R6083 IBIAS.n1 IBIAS.n0 9.3005
R6084 IBIAS.n24 IBIAS.n23 9.3005
R6085 IBIAS.n22 IBIAS.n21 9.3005
R6086 IBIAS.n20 IBIAS.n19 9.3005
R6087 IBIAS.n18 IBIAS.n17 9.3005
R6088 IBIAS.n16 IBIAS.n15 9.3005
R6089 IBIAS.n14 IBIAS.n13 9.3005
R6090 IBIAS.n12 IBIAS.n11 9.3005
R6091 IBIAS.n15 IBIAS.n5 8.28285
R6092 IBIAS.n17 IBIAS.n6 6.77697
R6093 IBIAS.n19 IBIAS.n7 5.27109
R6094 IBIAS IBIAS.n28 5.23142
R6095 IBIAS.n21 IBIAS.n8 3.76521
R6096 IBIAS.n26 IBIAS.t1 2.48621
R6097 IBIAS.n26 IBIAS.t2 2.48621
R6098 IBIAS.n10 IBIAS.n2 2.36936
R6099 IBIAS.n25 IBIAS.n24 2.25932
R6100 IBIAS.n10 IBIAS.n9 0.320353
R6101 IBIAS.n28 IBIAS.n0 0.196152
R6102 IBIAS.n23 IBIAS.n0 0.196152
R6103 IBIAS.n23 IBIAS.n22 0.196152
R6104 IBIAS.n22 IBIAS.n20 0.196152
R6105 IBIAS.n20 IBIAS.n18 0.196152
R6106 IBIAS.n18 IBIAS.n16 0.196152
R6107 IBIAS.n16 IBIAS.n14 0.196152
R6108 IBIAS.n14 IBIAS.n12 0.196152
R6109 IBIAS.n12 IBIAS.n10 0.196152
C0 VDD VOUT 9.72747f
C1 VP VOUT 0.48845f
C2 VP VN 5.95617f
C3 EN VOUT 0.69581f
C4 VOUT VN 0.15325f
C5 EN IBIAS 0.80192f
C6 C1 VDD 0.11857f
C7 C1 VOUT 57.8095f
C8 IBIAS VSS 1.96999f
C9 EN VSS 3.13615f
C10 VP VSS 5.19954f
C11 VN VSS 5.44205f
C12 VOUT VSS 20.47861f
C13 VDD VSS 14.74441f
C14 C1 VSS 33.84245f
C15 C1.t0 VSS 0.29149f
C16 C1.t1 VSS 28.5519f
C17 a_3758_2896.t6 VSS 0.03416f
C18 a_3758_2896.t3 VSS 0.03416f
C19 a_3758_2896.t4 VSS 0.03416f
C20 a_3758_2896.n0 VSS 0.11734f
C21 a_3758_2896.t0 VSS 0.03416f
C22 a_3758_2896.t10 VSS 0.03416f
C23 a_3758_2896.n1 VSS 0.10037f
C24 a_3758_2896.n2 VSS 0.75156f
C25 a_3758_2896.t9 VSS 0.03416f
C26 a_3758_2896.t8 VSS 0.03416f
C27 a_3758_2896.n3 VSS 0.10037f
C28 a_3758_2896.n4 VSS 0.39548f
C29 a_3758_2896.t2 VSS 0.03416f
C30 a_3758_2896.t1 VSS 0.03416f
C31 a_3758_2896.n5 VSS 0.10037f
C32 a_3758_2896.n6 VSS 0.39548f
C33 a_3758_2896.n7 VSS 0.01301f
C34 a_3758_2896.t14 VSS 0.12182f
C35 a_3758_2896.n9 VSS 0.01076f
C36 a_3758_2896.t13 VSS 0.79281f
C37 a_3758_2896.n16 VSS 1.50323f
C38 a_3758_2896.n17 VSS 0.21382f
C39 a_3758_2896.n19 VSS 0.01301f
C40 a_3758_2896.n21 VSS 0.01301f
C41 a_3758_2896.n23 VSS 0.01301f
C42 a_3758_2896.n25 VSS 0.01301f
C43 a_3758_2896.n27 VSS 0.01301f
C44 a_3758_2896.n29 VSS 0.01301f
C45 a_3758_2896.n30 VSS 0.01301f
C46 a_3758_2896.t12 VSS 0.07972f
C47 a_3758_2896.n33 VSS 0.17055f
C48 a_3758_2896.n35 VSS 0.36219f
C49 a_3758_2896.t5 VSS 0.03416f
C50 a_3758_2896.t7 VSS 0.03416f
C51 a_3758_2896.n36 VSS 0.10037f
C52 a_3758_2896.n37 VSS 0.64652f
C53 a_3758_2896.n38 VSS 0.33874f
C54 a_3758_2896.n39 VSS 0.10037f
C55 a_3758_2896.t11 VSS 0.03416f
C56 a_2479_9004.t3 VSS 0.02166f
C57 a_2479_9004.t1 VSS 0.02166f
C58 a_2479_9004.n0 VSS 0.04534f
C59 a_2479_9004.t23 VSS 0.09411f
C60 a_2479_9004.t2 VSS 0.09411f
C61 a_2479_9004.n1 VSS -0.15502f
C62 a_2479_9004.n2 VSS 0.2387f
C63 a_2479_9004.t24 VSS 0.09411f
C64 a_2479_9004.t0 VSS 0.09411f
C65 a_2479_9004.n3 VSS 0.24905f
C66 a_2479_9004.t6 VSS 0.09411f
C67 a_2479_9004.t21 VSS 0.09411f
C68 a_2479_9004.n4 VSS 0.24905f
C69 a_2479_9004.t4 VSS 0.09411f
C70 a_2479_9004.t16 VSS 0.1516f
C71 a_2479_9004.t15 VSS 0.1516f
C72 a_2479_9004.n5 VSS 0.84136f
C73 a_2479_9004.t20 VSS 0.1516f
C74 a_2479_9004.t19 VSS 0.1516f
C75 a_2479_9004.n6 VSS 0.62542f
C76 a_2479_9004.n7 VSS 3.09987f
C77 a_2479_9004.n8 VSS 0.02473f
C78 a_2479_9004.n9 VSS 0.01699f
C79 a_2479_9004.t17 VSS 0.1516f
C80 a_2479_9004.n10 VSS 0.02047f
C81 a_2479_9004.t10 VSS 0.08006f
C82 a_2479_9004.t8 VSS 1.50795f
C83 a_2479_9004.n17 VSS 2.88661f
C84 a_2479_9004.n18 VSS 0.40663f
C85 a_2479_9004.n19 VSS 0.01649f
C86 a_2479_9004.n20 VSS 0.02473f
C87 a_2479_9004.n22 VSS 0.02473f
C88 a_2479_9004.n24 VSS 0.02473f
C89 a_2479_9004.n26 VSS 0.02473f
C90 a_2479_9004.n28 VSS 0.02473f
C91 a_2479_9004.n30 VSS 0.02473f
C92 a_2479_9004.n31 VSS 0.02473f
C93 a_2479_9004.t9 VSS 0.1516f
C94 a_2479_9004.n34 VSS 0.32433f
C95 a_2479_9004.n35 VSS 0.01069f
C96 a_2479_9004.n36 VSS 0.38075f
C97 a_2479_9004.t14 VSS 0.1516f
C98 a_2479_9004.t13 VSS 0.1516f
C99 a_2479_9004.n37 VSS 0.61041f
C100 a_2479_9004.n38 VSS 1.4281f
C101 a_2479_9004.n39 VSS 0.02473f
C102 a_2479_9004.n40 VSS 0.01699f
C103 a_2479_9004.t12 VSS 0.23166f
C104 a_2479_9004.n41 VSS 0.02047f
C105 a_2479_9004.t11 VSS 1.50795f
C106 a_2479_9004.n48 VSS 2.88661f
C107 a_2479_9004.n49 VSS 0.40663f
C108 a_2479_9004.n50 VSS 0.01649f
C109 a_2479_9004.n51 VSS 0.02473f
C110 a_2479_9004.n53 VSS 0.02473f
C111 a_2479_9004.n55 VSS 0.02473f
C112 a_2479_9004.n57 VSS 0.02473f
C113 a_2479_9004.n59 VSS 0.02473f
C114 a_2479_9004.n61 VSS 0.02473f
C115 a_2479_9004.n62 VSS 0.02473f
C116 a_2479_9004.t18 VSS 0.1516f
C117 a_2479_9004.n65 VSS 0.32433f
C118 a_2479_9004.n66 VSS 0.01069f
C119 a_2479_9004.n67 VSS 0.19498f
C120 a_2479_9004.n68 VSS 0.36196f
C121 a_2479_9004.n69 VSS 1.87446f
C122 a_2479_9004.t22 VSS 0.09411f
C123 a_2479_9004.n70 VSS 0.94824f
C124 a_2479_9004.n71 VSS 0.2387f
C125 a_2479_9004.t5 VSS 0.02166f
C126 a_2479_9004.n72 VSS 0.04534f
C127 a_2479_9004.t7 VSS 0.02166f
C128 VN.t0 VSS 1.38469f
C129 VN.t1 VSS 1.38075f
C130 VN.n0 VSS 1.21869f
C131 VN.t4 VSS 1.38075f
C132 VN.n1 VSS 0.60854f
C133 VN.t5 VSS 1.38202f
C134 VN.n2 VSS 1.32742f
C135 VN.t7 VSS 1.38043f
C136 VN.t2 VSS 1.38365f
C137 VN.t6 VSS 1.38043f
C138 VN.n3 VSS 1.20405f
C139 VN.n4 VSS 0.57632f
C140 VN.t3 VSS 1.38021f
C141 VN.n5 VSS 0.59805f
C142 VN.n6 VSS 0.73649f
C143 a_2995_7336.t9 VSS 0.11279f
C144 a_2995_7336.t3 VSS 0.11279f
C145 a_2995_7336.t8 VSS 0.11279f
C146 a_2995_7336.n0 VSS 0.32268f
C147 a_2995_7336.t12 VSS 0.11279f
C148 a_2995_7336.t5 VSS 0.11279f
C149 a_2995_7336.n1 VSS 0.32268f
C150 a_2995_7336.t6 VSS 0.11279f
C151 a_2995_7336.t10 VSS 0.11279f
C152 a_2995_7336.n2 VSS 0.32272f
C153 a_2995_7336.n3 VSS 1.26812f
C154 a_2995_7336.t7 VSS 0.11279f
C155 a_2995_7336.t15 VSS 0.11279f
C156 a_2995_7336.n4 VSS 0.32268f
C157 a_2995_7336.t4 VSS 0.11279f
C158 a_2995_7336.t11 VSS 0.11279f
C159 a_2995_7336.n5 VSS 0.32272f
C160 a_2995_7336.n6 VSS 0.0184f
C161 a_2995_7336.n7 VSS 0.01264f
C162 a_2995_7336.t1 VSS 0.11279f
C163 a_2995_7336.n8 VSS 0.01523f
C164 a_2995_7336.t19 VSS 0.05957f
C165 a_2995_7336.t17 VSS 1.12173f
C166 a_2995_7336.n15 VSS 2.1269f
C167 a_2995_7336.n16 VSS 0.30254f
C168 a_2995_7336.n17 VSS 0.01227f
C169 a_2995_7336.n18 VSS 0.0184f
C170 a_2995_7336.n20 VSS 0.0184f
C171 a_2995_7336.n22 VSS 0.0184f
C172 a_2995_7336.n24 VSS 0.0184f
C173 a_2995_7336.n26 VSS 0.0184f
C174 a_2995_7336.n28 VSS 0.0184f
C175 a_2995_7336.n29 VSS 0.0184f
C176 a_2995_7336.t18 VSS 0.11279f
C177 a_2995_7336.n32 VSS 0.24131f
C178 a_2995_7336.n34 VSS 0.18922f
C179 a_2995_7336.t16 VSS 0.11279f
C180 a_2995_7336.t13 VSS 0.11279f
C181 a_2995_7336.n35 VSS 0.32268f
C182 a_2995_7336.t14 VSS 0.11279f
C183 a_2995_7336.t2 VSS 0.11279f
C184 a_2995_7336.n36 VSS 0.32272f
C185 a_2995_7336.n37 VSS 1.58502f
C186 a_2995_7336.n38 VSS 1.93909f
C187 a_2995_7336.n39 VSS 1.60509f
C188 a_2995_7336.n40 VSS 1.26814f
C189 a_2995_7336.n41 VSS 0.32269f
C190 a_2995_7336.t0 VSS 0.11279f
C191 VP.t7 VSS 1.38738f
C192 VP.t6 VSS 1.38343f
C193 VP.n0 VSS 1.22106f
C194 VP.t2 VSS 1.38343f
C195 VP.n1 VSS 0.60972f
C196 VP.t1 VSS 1.3847f
C197 VP.n2 VSS 1.27437f
C198 VP.t3 VSS 1.38633f
C199 VP.t5 VSS 1.38311f
C200 VP.n3 VSS 1.20639f
C201 VP.t4 VSS 1.38311f
C202 VP.n4 VSS 0.57744f
C203 VP.t0 VSS 1.38289f
C204 VP.n5 VSS 0.59921f
C205 VP.n6 VSS 0.717f
C206 a_4920_2896.t10 VSS 0.02015f
C207 a_4920_2896.t16 VSS 0.02015f
C208 a_4920_2896.n0 VSS 0.04651f
C209 a_4920_2896.t4 VSS 0.02015f
C210 a_4920_2896.t11 VSS 0.02015f
C211 a_4920_2896.n1 VSS 0.04651f
C212 a_4920_2896.t20 VSS 0.02015f
C213 a_4920_2896.t3 VSS 0.02015f
C214 a_4920_2896.n2 VSS 0.04651f
C215 a_4920_2896.t22 VSS 0.02015f
C216 a_4920_2896.t21 VSS 0.02015f
C217 a_4920_2896.n3 VSS 0.04651f
C218 a_4920_2896.t14 VSS 0.02015f
C219 a_4920_2896.t9 VSS 0.02015f
C220 a_4920_2896.n4 VSS 0.05823f
C221 a_4920_2896.n5 VSS 0.44309f
C222 a_4920_2896.n6 VSS 0.18382f
C223 a_4920_2896.n7 VSS 0.18382f
C224 a_4920_2896.n8 VSS 0.18382f
C225 a_4920_2896.t8 VSS 0.02015f
C226 a_4920_2896.t1 VSS 0.02015f
C227 a_4920_2896.n9 VSS 0.04759f
C228 a_4920_2896.t18 VSS 0.02015f
C229 a_4920_2896.t2 VSS 0.02015f
C230 a_4920_2896.n10 VSS 0.04759f
C231 a_4920_2896.t13 VSS 0.02015f
C232 a_4920_2896.t19 VSS 0.02015f
C233 a_4920_2896.n11 VSS 0.04759f
C234 a_4920_2896.t5 VSS 0.02015f
C235 a_4920_2896.t12 VSS 0.02015f
C236 a_4920_2896.n12 VSS 0.04759f
C237 a_4920_2896.t7 VSS 0.02015f
C238 a_4920_2896.t6 VSS 0.02015f
C239 a_4920_2896.n13 VSS 0.04759f
C240 a_4920_2896.t0 VSS 0.02015f
C241 a_4920_2896.t17 VSS 0.02015f
C242 a_4920_2896.n14 VSS 0.05955f
C243 a_4920_2896.n15 VSS 0.4586f
C244 a_4920_2896.n16 VSS 0.1917f
C245 a_4920_2896.n17 VSS 0.1917f
C246 a_4920_2896.n18 VSS 0.1917f
C247 a_4920_2896.n19 VSS 0.37064f
C248 a_4920_2896.t26 VSS 0.07185f
C249 a_4920_2896.t25 VSS 0.46761f
C250 a_4920_2896.n30 VSS 0.88664f
C251 a_4920_2896.n44 VSS 0.12612f
C252 a_4920_2896.t24 VSS 0.04702f
C253 a_4920_2896.n46 VSS 0.10059f
C254 a_4920_2896.n48 VSS 0.0652f
C255 a_4920_2896.n49 VSS 0.31283f
C256 a_4920_2896.n50 VSS 0.23403f
C257 a_4920_2896.t15 VSS 0.02015f
C258 a_4920_2896.n51 VSS 0.04651f
C259 a_4920_2896.t23 VSS 0.02015f
C260 a_2080_2896.t7 VSS 0.02936f
C261 a_2080_2896.t22 VSS 0.21364f
C262 a_2080_2896.t30 VSS 0.21316f
C263 a_2080_2896.n9 VSS 0.22163f
C264 a_2080_2896.t9 VSS 0.21316f
C265 a_2080_2896.n10 VSS 0.08384f
C266 a_2080_2896.t10 VSS 0.21316f
C267 a_2080_2896.n11 VSS 0.08384f
C268 a_2080_2896.t11 VSS 0.21316f
C269 a_2080_2896.n12 VSS 0.08384f
C270 a_2080_2896.t40 VSS 0.21316f
C271 a_2080_2896.n13 VSS 0.08384f
C272 a_2080_2896.t39 VSS 0.21316f
C273 a_2080_2896.n14 VSS 0.08384f
C274 a_2080_2896.t28 VSS 0.21316f
C275 a_2080_2896.n15 VSS 0.08384f
C276 a_2080_2896.t29 VSS 0.21316f
C277 a_2080_2896.n16 VSS 0.08384f
C278 a_2080_2896.t18 VSS 0.21316f
C279 a_2080_2896.n17 VSS 0.08384f
C280 a_2080_2896.t8 VSS 0.21316f
C281 a_2080_2896.n18 VSS 0.08384f
C282 a_2080_2896.t21 VSS 0.21316f
C283 a_2080_2896.n19 VSS 0.11277f
C284 a_2080_2896.t35 VSS 0.21356f
C285 a_2080_2896.t43 VSS 0.21238f
C286 a_2080_2896.t27 VSS 0.21229f
C287 a_2080_2896.n20 VSS 0.1205f
C288 a_2080_2896.n21 VSS 0.13801f
C289 a_2080_2896.t15 VSS 0.21238f
C290 a_2080_2896.t38 VSS 0.21229f
C291 a_2080_2896.n22 VSS 0.1205f
C292 a_2080_2896.n23 VSS 0.02104f
C293 a_2080_2896.t32 VSS 0.21238f
C294 a_2080_2896.t16 VSS 0.21229f
C295 a_2080_2896.n24 VSS 0.1205f
C296 a_2080_2896.n25 VSS 0.02104f
C297 a_2080_2896.t33 VSS 0.21238f
C298 a_2080_2896.t17 VSS 0.21229f
C299 a_2080_2896.n26 VSS 0.1205f
C300 a_2080_2896.n27 VSS 0.02104f
C301 a_2080_2896.t34 VSS 0.21238f
C302 a_2080_2896.t19 VSS 0.21229f
C303 a_2080_2896.n28 VSS 0.1205f
C304 a_2080_2896.n29 VSS 0.02104f
C305 a_2080_2896.n30 VSS 0.02104f
C306 a_2080_2896.t23 VSS 0.21238f
C307 a_2080_2896.n31 VSS 0.01136f
C308 a_2080_2896.t25 VSS 0.21238f
C309 a_2080_2896.n32 VSS 0.07247f
C310 a_2080_2896.n33 VSS 0.04758f
C311 a_2080_2896.t5 VSS 0.16153f
C312 a_2080_2896.t6 VSS 0.01258f
C313 a_2080_2896.t4 VSS 0.01258f
C314 a_2080_2896.n53 VSS 0.02517f
C315 a_2080_2896.n56 VSS 0.11181f
C316 a_2080_2896.t3 VSS 0.16153f
C317 a_2080_2896.n57 VSS 0.04758f
C318 a_2080_2896.n58 VSS 0.07247f
C319 a_2080_2896.n59 VSS 0.02104f
C320 a_2080_2896.t12 VSS 0.21238f
C321 a_2080_2896.t36 VSS 0.21229f
C322 a_2080_2896.n60 VSS 0.1205f
C323 a_2080_2896.n61 VSS 0.02104f
C324 a_2080_2896.t13 VSS 0.21238f
C325 a_2080_2896.t37 VSS 0.21229f
C326 a_2080_2896.n62 VSS 0.1205f
C327 a_2080_2896.n63 VSS 0.02104f
C328 a_2080_2896.t41 VSS 0.21238f
C329 a_2080_2896.t24 VSS 0.21229f
C330 a_2080_2896.n64 VSS 0.1205f
C331 a_2080_2896.n65 VSS 0.02104f
C332 a_2080_2896.t31 VSS 0.21238f
C333 a_2080_2896.t14 VSS 0.21229f
C334 a_2080_2896.n66 VSS 0.1205f
C335 a_2080_2896.n67 VSS 0.02104f
C336 a_2080_2896.t42 VSS 0.21238f
C337 a_2080_2896.t26 VSS 0.21229f
C338 a_2080_2896.n68 VSS 0.1205f
C339 a_2080_2896.n69 VSS 0.02104f
C340 a_2080_2896.t20 VSS 0.21316f
C341 a_2080_2896.n70 VSS 0.16653f
C342 a_2080_2896.n71 VSS 0.2988f
C343 a_2080_2896.n72 VSS 0.17452f
C344 a_2080_2896.t1 VSS 0.02936f
C345 a_2080_2896.n86 VSS 0.06282f
C346 a_2080_2896.n90 VSS 0.07876f
C347 a_2080_2896.t0 VSS 0.29202f
C348 a_2080_2896.n91 VSS 0.47059f
C349 a_2080_2896.n92 VSS 0.08427f
C350 a_2080_2896.t2 VSS 0.01433f
C351 VDD.t21 VSS 0.03732f
C352 VDD.t67 VSS 0.01297f
C353 VDD.n0 VSS 0.01159f
C354 VDD.t19 VSS 0.03446f
C355 VDD.n1 VSS 0.20128f
C356 VDD.n2 VSS 0.01757f
C357 VDD.n3 VSS 0.1863f
C358 VDD.n4 VSS 0.01757f
C359 VDD.n5 VSS 0.12582f
C360 VDD.n6 VSS 0.01757f
C361 VDD.n7 VSS 0.12582f
C362 VDD.n8 VSS 0.01757f
C363 VDD.n9 VSS 0.16729f
C364 VDD.n10 VSS 0.07089f
C365 VDD.n11 VSS 0.06005f
C366 VDD.n15 VSS 0.66468f
C367 VDD.n19 VSS 0.0133f
C368 VDD.t20 VSS 0.19482f
C369 VDD.n22 VSS 0.36385f
C370 VDD.n23 VSS 0.52429f
C371 VDD.n24 VSS 0.0133f
C372 VDD.n34 VSS 0.05235f
C373 VDD.n35 VSS 0.02031f
C374 VDD.t12 VSS 0.02945f
C375 VDD.n36 VSS 0.07599f
C376 VDD.n37 VSS 0.0254f
C377 VDD.t52 VSS 0.0345f
C378 VDD.n38 VSS 0.01947f
C379 VDD.n39 VSS 0.05962f
C380 VDD.t30 VSS 0.06761f
C381 VDD.n40 VSS 0.02497f
C382 VDD.n41 VSS 0.04085f
C383 VDD.t33 VSS 0.06759f
C384 VDD.n42 VSS 0.0254f
C385 VDD.n43 VSS 0.04085f
C386 VDD.t9 VSS 0.06763f
C387 VDD.n44 VSS 0.04504f
C388 VDD.n45 VSS 0.02031f
C389 VDD.n46 VSS 0.01652f
C390 VDD.t35 VSS 0.01586f
C391 VDD.n47 VSS 0.01652f
C392 VDD.t32 VSS 0.01586f
C393 VDD.n48 VSS 0.01654f
C394 VDD.t53 VSS 0.01586f
C395 VDD.n49 VSS 0.01654f
C396 VDD.n50 VSS 0.08188f
C397 VDD.n51 VSS 0.07908f
C398 VDD.n52 VSS 0.01757f
C399 VDD.n53 VSS 0.12582f
C400 VDD.n54 VSS 0.05235f
C401 VDD.t15 VSS 0.01586f
C402 VDD.n55 VSS 0.02497f
C403 VDD.n56 VSS 0.0254f
C404 VDD.t27 VSS 0.0345f
C405 VDD.t38 VSS 0.06763f
C406 VDD.t39 VSS 0.03738f
C407 VDD.n57 VSS 0.04504f
C408 VDD.n58 VSS 0.01652f
C409 VDD.n59 VSS 0.02031f
C410 VDD.n60 VSS 0.07599f
C411 VDD.n61 VSS 0.04085f
C412 VDD.t13 VSS 0.06759f
C413 VDD.n62 VSS 0.0254f
C414 VDD.n63 VSS 0.04085f
C415 VDD.t49 VSS 0.06761f
C416 VDD.n64 VSS 0.05962f
C417 VDD.n65 VSS 0.01947f
C418 VDD.n66 VSS 0.02031f
C419 VDD.n67 VSS 0.01652f
C420 VDD.t51 VSS 0.01586f
C421 VDD.n68 VSS 0.01654f
C422 VDD.t29 VSS 0.01586f
C423 VDD.n69 VSS 0.01654f
C424 VDD.n70 VSS 0.08188f
C425 VDD.n71 VSS 0.11722f
C426 VDD.n72 VSS 0.05197f
C427 VDD.n100 VSS 0.06005f
C428 VDD.n115 VSS 0.01366f
C429 VDD.n116 VSS 0.01366f
C430 VDD.n117 VSS 0.0133f
C431 VDD.t14 VSS 0.19482f
C432 VDD.n123 VSS 0.37531f
C433 VDD.t28 VSS 0.19482f
C434 VDD.n130 VSS 0.38677f
C435 VDD.t0 VSS 0.19482f
C436 VDD.t7 VSS 0.19482f
C437 VDD.n140 VSS 0.38677f
C438 VDD.t17 VSS 0.19482f
C439 VDD.n147 VSS 0.37531f
C440 VDD.t34 VSS 0.19482f
C441 VDD.n152 VSS 0.0133f
C442 VDD.n153 VSS 0.0133f
C443 VDD.n154 VSS 0.36385f
C444 VDD.n156 VSS 0.0133f
C445 VDD.n168 VSS 0.01366f
C446 VDD.n172 VSS 0.03112f
C447 VDD.n176 VSS 0.02339f
C448 VDD.n204 VSS 0.0133f
C449 VDD.n205 VSS 0.01366f
C450 VDD.n240 VSS 0.09173f
C451 VDD.n241 VSS 0.0323f
C452 VDD.n252 VSS 0.09407f
C453 VDD.n255 VSS 0.01366f
C454 VDD.n256 VSS 0.01366f
C455 VDD.n258 VSS 0.66468f
C456 VDD.n259 VSS 0.52429f
C457 VDD.t10 VSS 0.19482f
C458 VDD.n260 VSS 0.22634f
C459 VDD.n266 VSS 0.2206f
C460 VDD.n267 VSS 0.36958f
C461 VDD.t31 VSS 0.19482f
C462 VDD.n268 VSS 0.21487f
C463 VDD.n274 VSS 0.20915f
C464 VDD.n275 VSS 0.38104f
C465 VDD.t2 VSS 0.19482f
C466 VDD.n276 VSS 0.20341f
C467 VDD.n282 VSS 0.19769f
C468 VDD.n283 VSS 0.38964f
C469 VDD.n284 VSS 0.19769f
C470 VDD.n290 VSS 0.20341f
C471 VDD.t5 VSS 0.19482f
C472 VDD.n291 VSS 0.38104f
C473 VDD.n292 VSS 0.20915f
C474 VDD.n298 VSS 0.21487f
C475 VDD.t50 VSS 0.19482f
C476 VDD.n299 VSS 0.36958f
C477 VDD.n300 VSS 0.2206f
C478 VDD.n306 VSS 0.22634f
C479 VDD.n309 VSS 0.0133f
C480 VDD.n310 VSS 0.01366f
C481 VDD.n311 VSS 0.01366f
C482 VDD.n324 VSS 0.05234f
C483 VDD.n325 VSS 0.05235f
C484 VDD.t26 VSS 0.01586f
C485 VDD.n326 VSS 0.01947f
C486 VDD.n327 VSS 0.07599f
C487 VDD.n328 VSS 0.04085f
C488 VDD.t47 VSS 0.06763f
C489 VDD.t48 VSS 0.03738f
C490 VDD.n329 VSS 0.01652f
C491 VDD.n330 VSS 0.02031f
C492 VDD.n331 VSS 0.04504f
C493 VDD.n332 VSS 0.0254f
C494 VDD.t25 VSS 0.06759f
C495 VDD.n333 VSS 0.0254f
C496 VDD.t36 VSS 0.0345f
C497 VDD.n334 VSS 0.05962f
C498 VDD.t54 VSS 0.06761f
C499 VDD.n335 VSS 0.04085f
C500 VDD.n336 VSS 0.02497f
C501 VDD.n337 VSS 0.02031f
C502 VDD.n338 VSS 0.01652f
C503 VDD.t55 VSS 0.01586f
C504 VDD.n339 VSS 0.01654f
C505 VDD.t37 VSS 0.01586f
C506 VDD.n340 VSS 0.01654f
C507 VDD.n341 VSS 0.08188f
C508 VDD.n342 VSS 0.11777f
C509 VDD.n343 VSS 0.01757f
C510 VDD.n344 VSS 0.12582f
C511 VDD.n345 VSS 0.05235f
C512 VDD.n346 VSS 0.02031f
C513 VDD.n347 VSS 0.04504f
C514 VDD.n348 VSS 0.02497f
C515 VDD.t24 VSS 0.02945f
C516 VDD.n349 VSS 0.04085f
C517 VDD.t16 VSS 0.0345f
C518 VDD.t40 VSS 0.06761f
C519 VDD.n350 VSS 0.05962f
C520 VDD.n351 VSS 0.01947f
C521 VDD.n352 VSS 0.0254f
C522 VDD.t45 VSS 0.06759f
C523 VDD.n353 VSS 0.0254f
C524 VDD.t22 VSS 0.06763f
C525 VDD.n354 VSS 0.04085f
C526 VDD.n355 VSS 0.07599f
C527 VDD.n356 VSS 0.02031f
C528 VDD.n357 VSS 0.01652f
C529 VDD.t46 VSS 0.01586f
C530 VDD.n358 VSS 0.01652f
C531 VDD.t41 VSS 0.01586f
C532 VDD.n359 VSS 0.01654f
C533 VDD.t18 VSS 0.01586f
C534 VDD.n360 VSS 0.01654f
C535 VDD.n361 VSS 0.08188f
C536 VDD.n362 VSS 0.09929f
C537 VDD.n363 VSS 0.01815f
C538 VDD.n364 VSS 0.01757f
C539 VDD.n365 VSS 0.32102f
C540 VDD.n366 VSS 0.01757f
C541 VDD.n367 VSS 0.12582f
C542 VDD.n368 VSS 0.01757f
C543 VDD.n369 VSS 0.12582f
C544 VDD.t44 VSS 0.02939f
C545 VDD.n370 VSS 0.01654f
C546 VDD.n371 VSS 0.1123f
C547 VDD.t42 VSS 0.03446f
C548 VDD.n372 VSS 0.07395f
C549 VDD.n373 VSS 0.10279f
C550 VDD.n374 VSS 0.41359f
C551 VDD.n375 VSS 0.26431f
C552 VDD.n376 VSS 0.19985f
C553 VOUT.n0 VSS 0.01561f
C554 VOUT.n1 VSS 0.01513f
C555 VOUT.n2 VSS 0.2765f
C556 VOUT.n3 VSS 0.01513f
C557 VOUT.n4 VSS 0.11605f
C558 VOUT.n5 VSS 0.01513f
C559 VOUT.n6 VSS 0.11605f
C560 VOUT.n7 VSS 0.03194f
C561 VOUT.n8 VSS 0.03838f
C562 VOUT.t8 VSS 0.05763f
C563 VOUT.t10 VSS 0.02509f
C564 VOUT.n9 VSS 0.01408f
C565 VOUT.t5 VSS 0.01351f
C566 VOUT.n10 VSS 0.01408f
C567 VOUT.n11 VSS 0.01731f
C568 VOUT.n12 VSS 0.06898f
C569 VOUT.n13 VSS 0.0566f
C570 VOUT.t4 VSS 0.05761f
C571 VOUT.n14 VSS 0.02164f
C572 VOUT.n15 VSS 0.04613f
C573 VOUT.n16 VSS 0.10296f
C574 VOUT.t0 VSS 0.04729f
C575 VOUT.t13 VSS 0.02497f
C576 VOUT.t11 VSS 0.47028f
C577 VOUT.n26 VSS 0.89169f
C578 VOUT.n27 VSS 0.12684f
C579 VOUT.t12 VSS 0.04729f
C580 VOUT.n43 VSS 0.10117f
C581 VOUT.n45 VSS 0.44202f
C582 VOUT.n46 VSS 0.66145f
C583 VOUT.n48 VSS 0.01789f
C584 VOUT.t1 VSS 66.8769f
C585 VOUT.n49 VSS 0.03885f
C586 VOUT.n50 VSS 0.03489f
C587 VOUT.n51 VSS 1.16187f
C588 VOUT.n52 VSS 0.02957f
C589 VOUT.n53 VSS 0.02031f
C590 VOUT.n54 VSS 0.02041f
C591 VOUT.n55 VSS 0.06898f
C592 VOUT.t3 VSS 0.03185f
C593 VOUT.t6 VSS 0.05761f
C594 VOUT.n56 VSS 0.0566f
C595 VOUT.t2 VSS 0.05763f
C596 VOUT.n57 VSS 0.03838f
C597 VOUT.n58 VSS 0.01731f
C598 VOUT.n59 VSS 0.01408f
C599 VOUT.t7 VSS 0.01351f
C600 VOUT.n60 VSS 0.01408f
C601 VOUT.n61 VSS 0.0334f
C602 VOUT.n62 VSS 0.06133f
C603 VOUT.n63 VSS 0.01513f
C604 VOUT.n64 VSS 0.18517f
C605 VOUT.n65 VSS 0.01513f
C606 VOUT.n66 VSS 0.11605f
C607 VOUT.n67 VSS 0.01513f
C608 VOUT.n68 VSS 0.11605f
C609 VOUT.n69 VSS 0.01513f
C610 VOUT.n70 VSS 0.16056f
C611 VOUT.n71 VSS 0.27023f
C612 VOUT.n72 VSS 0.3823f
C613 a_2479_7336.t9 VSS 0.0167f
C614 a_2479_7336.t31 VSS 0.07266f
C615 a_2479_7336.t22 VSS 0.07257f
C616 a_2479_7336.n0 VSS 0.13473f
C617 a_2479_7336.t24 VSS 0.07257f
C618 a_2479_7336.n1 VSS 0.06264f
C619 a_2479_7336.n2 VSS 0.01907f
C620 a_2479_7336.n3 VSS 0.0131f
C621 a_2479_7336.t14 VSS 0.17862f
C622 a_2479_7336.n11 VSS 0.01271f
C623 a_2479_7336.t13 VSS 1.16271f
C624 a_2479_7336.n12 VSS 2.22574f
C625 a_2479_7336.n14 VSS 0.01907f
C626 a_2479_7336.n16 VSS 0.01907f
C627 a_2479_7336.n18 VSS 0.01907f
C628 a_2479_7336.n20 VSS 0.01907f
C629 a_2479_7336.n22 VSS 0.01907f
C630 a_2479_7336.n24 VSS 0.01907f
C631 a_2479_7336.n25 VSS 0.01907f
C632 a_2479_7336.n26 VSS 0.31354f
C633 a_2479_7336.n27 VSS 0.01578f
C634 a_2479_7336.t7 VSS 0.11689f
C635 a_2479_7336.n28 VSS 0.25008f
C636 a_2479_7336.n30 VSS 0.29352f
C637 a_2479_7336.t16 VSS 0.11689f
C638 a_2479_7336.t6 VSS 0.11689f
C639 a_2479_7336.n31 VSS 0.47063f
C640 a_2479_7336.n32 VSS 1.10123f
C641 a_2479_7336.n33 VSS 0.01907f
C642 a_2479_7336.n34 VSS 0.0131f
C643 a_2479_7336.t15 VSS 0.11689f
C644 a_2479_7336.n42 VSS 0.01271f
C645 a_2479_7336.t12 VSS 0.06173f
C646 a_2479_7336.t10 VSS 1.16271f
C647 a_2479_7336.n43 VSS 2.22574f
C648 a_2479_7336.n45 VSS 0.01907f
C649 a_2479_7336.n47 VSS 0.01907f
C650 a_2479_7336.n49 VSS 0.01907f
C651 a_2479_7336.n51 VSS 0.01907f
C652 a_2479_7336.n53 VSS 0.01907f
C653 a_2479_7336.n55 VSS 0.01907f
C654 a_2479_7336.n56 VSS 0.01907f
C655 a_2479_7336.n57 VSS 0.31354f
C656 a_2479_7336.n58 VSS 0.01578f
C657 a_2479_7336.t11 VSS 0.11689f
C658 a_2479_7336.n59 VSS 0.25008f
C659 a_2479_7336.n61 VSS 0.15034f
C660 a_2479_7336.n62 VSS 1.04669f
C661 a_2479_7336.t5 VSS 0.11689f
C662 a_2479_7336.t4 VSS 0.11689f
C663 a_2479_7336.n63 VSS 0.48226f
C664 a_2479_7336.n64 VSS 1.6235f
C665 a_2479_7336.t3 VSS 0.11689f
C666 a_2479_7336.t2 VSS 0.11689f
C667 a_2479_7336.n65 VSS 0.48226f
C668 a_2479_7336.n66 VSS 1.41356f
C669 a_2479_7336.t17 VSS 0.0167f
C670 a_2479_7336.t1 VSS 0.0167f
C671 a_2479_7336.n67 VSS 0.03522f
C672 a_2479_7336.t19 VSS 0.07266f
C673 a_2479_7336.t28 VSS 0.07257f
C674 a_2479_7336.n68 VSS 0.13473f
C675 a_2479_7336.t35 VSS 0.07257f
C676 a_2479_7336.n69 VSS 0.06264f
C677 a_2479_7336.n70 VSS 0.16286f
C678 a_2479_7336.t32 VSS 0.07257f
C679 a_2479_7336.n71 VSS 0.06264f
C680 a_2479_7336.t26 VSS 0.07257f
C681 a_2479_7336.n72 VSS 0.07178f
C682 a_2479_7336.t23 VSS 0.07257f
C683 a_2479_7336.n73 VSS 0.07178f
C684 a_2479_7336.t20 VSS 0.07257f
C685 a_2479_7336.n74 VSS 0.07178f
C686 a_2479_7336.t30 VSS 0.07257f
C687 a_2479_7336.n75 VSS 0.07178f
C688 a_2479_7336.t25 VSS 0.07257f
C689 a_2479_7336.n76 VSS 0.12224f
C690 a_2479_7336.t8 VSS 0.718f
C691 a_2479_7336.n77 VSS 5.01875f
C692 a_2479_7336.n78 VSS 2.41673f
C693 a_2479_7336.t34 VSS 0.07257f
C694 a_2479_7336.n79 VSS 0.1168f
C695 a_2479_7336.t21 VSS 0.07257f
C696 a_2479_7336.n80 VSS 0.07178f
C697 a_2479_7336.t29 VSS 0.07257f
C698 a_2479_7336.n81 VSS 0.07178f
C699 a_2479_7336.t18 VSS 0.07257f
C700 a_2479_7336.n82 VSS 0.07178f
C701 a_2479_7336.t33 VSS 0.07257f
C702 a_2479_7336.n83 VSS 0.07178f
C703 a_2479_7336.t27 VSS 0.07257f
C704 a_2479_7336.n84 VSS 0.06264f
C705 a_2479_7336.n85 VSS 0.16286f
C706 a_2479_7336.n86 VSS 0.03522f
C707 a_2479_7336.t0 VSS 0.0167f
.ends

