* NGSPICE file created from two_stage_op_amp.ext - technology: sky130A

.subckt two_stage_op_amp IBIAS EN VOUT VN VP VDD VSS
X0 VDD.t31 a_2479_7336.t18 VOUT.t0 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X1 VSS.t172 VSS.t171 VSS.t172 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X2 VSS.t170 VSS.t169 VSS.t170 VSS.t42 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X3 VDD.t30 a_2479_7336.t19 VOUT.t14 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X4 VDD.t76 VDD.t75 VDD.t76 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X5 VSS.t168 VSS.t167 a_4920_2896.t25 VSS.t84 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X6 VSS.t160 VSS.t159 a_4920_2896.t24 VSS.t81 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X7 a_2479_7336.t11 a_2479_7336.t10 a_2479_7336.t11 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X8 VSS.t166 VSS.t165 VSS.t166 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X9 VDD.t74 VDD.t73 VDD.t74 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X10 VDD.t29 a_2479_7336.t20 VOUT.t2 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X11 VDD.t28 a_2479_7336.t21 VOUT.t13 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X12 a_4920_2896.t23 VSS.t163 VSS.t164 VSS.t78 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X13 a_2479_7336.t9 a_2479_7336.t7 a_2479_7336.t8 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X14 a_2479_7336.t3 VP.t0 a_2995_7336.t8 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X15 VSS.t162 VSS.t161 a_4920_2896.t22 VSS.t75 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X16 VSS.t158 VSS.t157 VSS.t158 VSS.t72 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X17 a_2995_7336.t14 VN.t0 a_2479_9004.t20 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X18 VDD.t26 a_2479_7336.t22 VOUT.t9 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X19 a_2479_9004.t19 VN.t1 a_2995_7336.t19 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X20 VSS.t156 VSS.t155 VSS.t156 VSS.t66 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X21 a_2479_9004.t4 a_2479_9004.t3 a_2479_9004.t4 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X22 VSS.t154 VSS.t153 VSS.t154 VSS.t69 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X23 a_4920_2896.t21 VSS.t151 VSS.t152 VSS.t63 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X24 a_2479_9004.t2 a_2479_9004.t0 a_2479_9004.t1 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X25 a_2479_9004.t18 VN.t2 a_2995_7336.t15 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X26 VSS.t150 VSS.t149 a_4920_2896.t20 VSS.t57 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X27 VOUT.t15 a_2479_7336.t23 VDD.t24 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X28 VSS.t148 VSS.t147 VSS.t148 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X29 VDD.t72 VDD.t71 VDD.t72 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X30 a_2995_7336.t7 VP.t1 a_2479_7336.t4 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X31 VSS.t146 VSS.t145 VSS.t146 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X32 a_3758_2896.t13 VSS.t143 VSS.t144 VSS.t84 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X33 a_4920_2896.t19 VSS.t117 VSS.t118 VSS.t54 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X34 a_2479_7336.t2 VP.t2 a_2995_7336.t6 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X35 a_3758_2896.t12 VSS.t133 VSS.t134 VSS.t81 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X36 VOUT.t4 a_2479_7336.t24 VDD.t23 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X37 VSS.t142 VSS.t141 a_3758_2896.t11 VSS.t78 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X38 a_4920_2896.t1 a_4920_2896.t0 a_4920_2896.t1 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X39 a_4920_2896.t18 VSS.t139 VSS.t140 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X40 a_3758_2896.t10 VSS.t137 VSS.t138 VSS.t75 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X41 a_3758_2896.t9 VSS.t135 VSS.t136 VSS.t72 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X42 a_4920_2896.t26 EN.t0 VOUT.t33 VSS.t177 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X43 a_2995_7336.t5 VP.t3 a_2479_7336.t6 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X44 VDD.t34 a_2479_9004.t11 a_2479_9004.t12 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X45 VOUT.t31 VOUT.t29 VOUT.t30 VSS.t173 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X46 a_4920_2896.t17 VSS.t131 VSS.t132 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X47 VDD.t70 VDD.t69 VDD.t70 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X48 VSS.t17 VSS.t15 a_4920_2896.t16 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X49 VDD.t68 VDD.t67 VDD.t68 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X50 VSS.t130 VSS.t129 VSS.t130 VSS.t111 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X51 VDD.t22 a_2479_7336.t25 VOUT.t10 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X52 VSS.t128 VSS.t126 VSS.t127 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X53 VSS.t116 VSS.t115 VSS.t116 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X54 VOUT.t28 VOUT.t26 VOUT.t27 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X55 VSS.t125 VSS.t124 a_4920_2896.t15 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X56 VOUT.t25 VOUT.t24 VOUT.t25 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X57 a_2995_7336.t17 VN.t3 a_2479_9004.t17 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X58 VDD.t20 a_2479_7336.t26 VOUT.t7 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X59 VSS.t123 VSS.t121 VSS.t122 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X60 VDD.t66 VDD.t64 VDD.t65 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X61 a_2479_9004.t10 a_2479_9004.t9 VDD.t4 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X62 VOUT.t18 VOUT.t19 sky130_fd_pr__cap_mim_m3_1 l=25.5 w=25.5
X63 VDD.t19 a_2479_7336.t27 VOUT.t17 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X64 VSS.t120 VSS.t119 a_3758_2896.t8 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X65 a_4920_2896.t14 VSS.t113 VSS.t114 VSS.t42 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X66 VSS.t112 VSS.t110 VSS.t112 VSS.t111 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X67 VOUT.t16 a_2479_7336.t28 VDD.t17 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X68 VDD.t3 a_2479_9004.t21 a_2479_7336.t1 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X69 VDD.t63 VDD.t62 VDD.t63 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X70 VSS.t109 VSS.t108 VSS.t109 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X71 VDD.t61 VDD.t60 VDD.t61 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X72 VOUT.t5 a_2479_7336.t29 VDD.t16 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X73 VSS.t14 VSS.t12 a_3758_2896.t7 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X74 VSS.t107 VSS.t106 VSS.t107 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X75 VDD.t59 VDD.t58 VDD.t59 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X76 VSS.t48 VSS.t47 VSS.t48 VSS.t45 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X77 VDD.t57 VDD.t56 VDD.t57 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X78 a_3758_2896.t6 VSS.t104 VSS.t105 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X79 VSS.t103 VSS.t102 VSS.t103 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X80 VSS.t101 VSS.t100 VSS.t101 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X81 VSS.t99 VSS.t98 VSS.t99 VSS.t66 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X82 a_2995_7336.t4 VP.t4 a_2479_7336.t15 VSS.t111 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X83 VSS.t97 VSS.t96 VSS.t97 VSS.t69 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X84 a_4920_2896.t13 VSS.t94 VSS.t95 VSS.t63 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X85 a_2479_7336.t12 VP.t5 a_2995_7336.t3 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X86 VSS.t93 VSS.t90 VSS.t92 VSS.t91 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X87 a_2479_7336.t0 a_2479_9004.t22 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X88 VSS.t89 VSS.t88 a_4920_2896.t12 VSS.t57 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X89 a_2995_7336.t18 VN.t4 a_2479_9004.t16 VSS.t45 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X90 VOUT.t11 a_2479_7336.t30 VDD.t14 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X91 a_4920_2896.t11 VSS.t86 VSS.t87 VSS.t54 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X92 a_2479_9004.t15 VN.t5 a_2995_7336.t13 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X93 VDD.t37 a_2479_9004.t23 a_2479_7336.t17 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X94 VDD.t55 VDD.t54 VDD.t55 VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X95 VSS.t85 VSS.t83 a_4920_2896.t10 VSS.t84 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X96 VOUT.t8 a_2479_7336.t31 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X97 VSS.t82 VSS.t80 a_4920_2896.t9 VSS.t81 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X98 a_2995_7336.t12 VN.t6 a_2479_9004.t14 VSS.t111 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X99 VDD.t53 VDD.t52 VDD.t53 VDD.t25 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X100 a_4920_2896.t8 VSS.t77 VSS.t79 VSS.t78 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X101 a_2479_9004.t13 VN.t7 a_2995_7336.t0 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X102 VSS.t76 VSS.t74 a_4920_2896.t7 VSS.t75 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X103 VSS.t73 VSS.t71 VSS.t73 VSS.t72 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X104 a_2995_7336.t2 VP.t6 a_2479_7336.t13 VSS.t45 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X105 a_2479_7336.t5 VP.t7 a_2995_7336.t1 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X106 VSS.t67 VSS.t65 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X107 VSS.t70 VSS.t68 a_3758_2896.t5 VSS.t69 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X108 VSS.t64 VSS.t62 a_3758_2896.t4 VSS.t63 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X109 VSS.t61 VSS.t59 VSS.t60 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X110 a_3758_2896.t3 VSS.t56 VSS.t58 VSS.t57 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X111 VDD.t6 a_2479_9004.t7 a_2479_9004.t8 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X112 VSS.t55 VSS.t53 a_3758_2896.t2 VSS.t54 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X113 IBIAS.t2 IBIAS.t1 IBIAS.t2 VSS.t176 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X114 VSS.t52 VSS.t51 VSS.t52 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X115 VDD.t51 VDD.t50 VDD.t51 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X116 VSS.t50 VSS.t49 a_4920_2896.t6 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X117 VDD.t49 VDD.t47 VDD.t48 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X118 IBIAS.t0 EN.t1 VSS.t180 VSS.t179 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X119 VSS.t46 VSS.t44 VSS.t46 VSS.t45 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X120 a_2479_7336.t16 a_2479_9004.t24 VDD.t35 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X121 a_4920_2896.t5 VSS.t41 VSS.t43 VSS.t42 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X122 a_4920_2896.t4 VSS.t38 VSS.t40 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X123 VOUT.t12 a_2479_7336.t32 VDD.t11 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X124 VDD.t46 VDD.t45 VDD.t46 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X125 VDD.t44 VDD.t43 VDD.t44 VDD.t15 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X126 a_3758_2896.t1 a_3758_2896.t0 a_3758_2896.t1 VSS.t174 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X127 VOUT.t6 a_2479_7336.t33 VDD.t10 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X128 VOUT.t23 VOUT.t22 VOUT.t23 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X129 a_4920_2896.t3 VSS.t36 VSS.t37 VSS.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X130 a_3758_2896.t14 EN.t2 a_2995_7336.t16 VSS.t178 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=1
X131 VSS.t35 VSS.t34 a_4920_2896.t2 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=1
X132 VOUT.t21 VOUT.t20 VOUT.t21 VDD.t32 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X133 VOUT.t1 a_2479_7336.t34 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X134 VSS.t33 VSS.t30 VSS.t32 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=0.87 pd=6.58 as=0 ps=0 w=3 l=1
X135 a_2995_7336.t11 a_2995_7336.t9 a_2995_7336.t10 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X136 VDD.t42 VDD.t41 VDD.t42 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0 ps=0 w=1 l=0.4
X137 VSS.t29 VSS.t28 VSS.t29 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X138 VDD.t40 VDD.t38 VDD.t39 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.4
X139 a_2479_7336.t14 VOUT.t32 VSS.t175 sky130_fd_pr__res_xhigh_po_1p41 l=14
X140 VSS.t27 VSS.t25 VSS.t27 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=0.435 pd=3.29 as=0 ps=0 w=3 l=1
X141 VSS.t24 VSS.t22 VSS.t23 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=2.03 pd=14.58 as=0 ps=0 w=7 l=1
X142 VSS.t21 VSS.t20 VSS.t21 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X143 VDD.t7 a_2479_7336.t35 VOUT.t3 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X144 VSS.t19 VSS.t18 VSS.t19 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
X145 a_2479_9004.t6 a_2479_9004.t5 VDD.t36 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.29 as=0.145 ps=1.29 w=1 l=0.4
X146 VSS.t11 VSS.t10 VSS.t11 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.015 pd=7.29 as=0 ps=0 w=7 l=1
C0 VOUT VN 0.15325f
C1 VOUT VP 0.38099f
C2 VOUT EN 0.69581f
C3 VDD VOUT 9.68294f
C4 VN VP 5.95617f
C5 IBIAS EN 0.80152f
R0 a_2479_7336.n83 a_2479_7336.t19 260.486
R1 a_2479_7336.n66 a_2479_7336.t31 260.486
R2 a_2479_7336.n83 a_2479_7336.t28 260.111
R3 a_2479_7336.n84 a_2479_7336.t35 260.111
R4 a_2479_7336.n82 a_2479_7336.t32 260.111
R5 a_2479_7336.n81 a_2479_7336.t26 260.111
R6 a_2479_7336.n80 a_2479_7336.t23 260.111
R7 a_2479_7336.n79 a_2479_7336.t20 260.111
R8 a_2479_7336.n78 a_2479_7336.t30 260.111
R9 a_2479_7336.n77 a_2479_7336.t25 260.111
R10 a_2479_7336.n74 a_2479_7336.t34 260.111
R11 a_2479_7336.n73 a_2479_7336.t21 260.111
R12 a_2479_7336.n72 a_2479_7336.t29 260.111
R13 a_2479_7336.n71 a_2479_7336.t18 260.111
R14 a_2479_7336.n70 a_2479_7336.t33 260.111
R15 a_2479_7336.n69 a_2479_7336.t27 260.111
R16 a_2479_7336.n67 a_2479_7336.t24 260.111
R17 a_2479_7336.n66 a_2479_7336.t22 260.111
R18 a_2479_7336.n68 a_2479_7336.n65 203.843
R19 a_2479_7336.n86 a_2479_7336.n85 203.841
R20 a_2479_7336.n57 a_2479_7336.n39 185
R21 a_2479_7336.n57 a_2479_7336.n38 185
R22 a_2479_7336.n57 a_2479_7336.n37 185
R23 a_2479_7336.n57 a_2479_7336.n36 185
R24 a_2479_7336.n57 a_2479_7336.n35 185
R25 a_2479_7336.n57 a_2479_7336.n34 185
R26 a_2479_7336.n57 a_2479_7336.n33 185
R27 a_2479_7336.n26 a_2479_7336.n8 185
R28 a_2479_7336.n26 a_2479_7336.n7 185
R29 a_2479_7336.n26 a_2479_7336.n6 185
R30 a_2479_7336.n26 a_2479_7336.n5 185
R31 a_2479_7336.n26 a_2479_7336.n4 185
R32 a_2479_7336.n26 a_2479_7336.n3 185
R33 a_2479_7336.n26 a_2479_7336.n2 185
R34 a_2479_7336.n41 a_2479_7336.t7 130.75
R35 a_2479_7336.n10 a_2479_7336.t10 130.75
R36 a_2479_7336.n41 a_2479_7336.t9 91.3557
R37 a_2479_7336.n10 a_2479_7336.t11 91.3557
R38 a_2479_7336.n58 a_2479_7336.n57 86.5152
R39 a_2479_7336.n27 a_2479_7336.n26 86.5152
R40 a_2479_7336.n56 a_2479_7336.n40 30.3012
R41 a_2479_7336.n25 a_2479_7336.n9 30.3012
R42 a_2479_7336.n65 a_2479_7336.t17 28.5655
R43 a_2479_7336.n65 a_2479_7336.t16 28.5655
R44 a_2479_7336.n86 a_2479_7336.t1 28.5655
R45 a_2479_7336.t0 a_2479_7336.n86 28.5655
R46 a_2479_7336.n33 a_2479_7336.n32 24.8476
R47 a_2479_7336.n2 a_2479_7336.n1 24.8476
R48 a_2479_7336.n42 a_2479_7336.n34 23.3417
R49 a_2479_7336.n11 a_2479_7336.n3 23.3417
R50 a_2479_7336.n59 a_2479_7336.n58 22.0256
R51 a_2479_7336.n28 a_2479_7336.n27 22.0256
R52 a_2479_7336.n44 a_2479_7336.n35 21.8358
R53 a_2479_7336.n13 a_2479_7336.n4 21.8358
R54 a_2479_7336.n46 a_2479_7336.n36 20.3299
R55 a_2479_7336.n15 a_2479_7336.n5 20.3299
R56 a_2479_7336.n48 a_2479_7336.n37 18.824
R57 a_2479_7336.n17 a_2479_7336.n6 18.824
R58 a_2479_7336.n50 a_2479_7336.n38 17.3181
R59 a_2479_7336.n19 a_2479_7336.n7 17.3181
R60 a_2479_7336.n57 a_2479_7336.n56 16.3559
R61 a_2479_7336.n26 a_2479_7336.n25 16.3559
R62 a_2479_7336.n52 a_2479_7336.n39 15.8123
R63 a_2479_7336.n21 a_2479_7336.n8 15.8123
R64 a_2479_7336.n62 a_2479_7336.n61 14.6052
R65 a_2479_7336.n64 a_2479_7336.n63 14.6052
R66 a_2479_7336.n30 a_2479_7336.n29 14.377
R67 a_2479_7336.n58 a_2479_7336.n32 12.7256
R68 a_2479_7336.n27 a_2479_7336.n1 12.7256
R69 a_2479_7336.n62 a_2479_7336.n60 11.5586
R70 a_2479_7336.n40 a_2479_7336.n39 11.2946
R71 a_2479_7336.n9 a_2479_7336.n8 11.2946
R72 a_2479_7336.n52 a_2479_7336.n38 9.78874
R73 a_2479_7336.n21 a_2479_7336.n7 9.78874
R74 a_2479_7336.n32 a_2479_7336.n31 9.3005
R75 a_2479_7336.n43 a_2479_7336.n42 9.3005
R76 a_2479_7336.n45 a_2479_7336.n44 9.3005
R77 a_2479_7336.n47 a_2479_7336.n46 9.3005
R78 a_2479_7336.n49 a_2479_7336.n48 9.3005
R79 a_2479_7336.n51 a_2479_7336.n50 9.3005
R80 a_2479_7336.n53 a_2479_7336.n52 9.3005
R81 a_2479_7336.n54 a_2479_7336.n40 9.3005
R82 a_2479_7336.n1 a_2479_7336.n0 9.3005
R83 a_2479_7336.n12 a_2479_7336.n11 9.3005
R84 a_2479_7336.n14 a_2479_7336.n13 9.3005
R85 a_2479_7336.n16 a_2479_7336.n15 9.3005
R86 a_2479_7336.n18 a_2479_7336.n17 9.3005
R87 a_2479_7336.n20 a_2479_7336.n19 9.3005
R88 a_2479_7336.n22 a_2479_7336.n21 9.3005
R89 a_2479_7336.n23 a_2479_7336.n9 9.3005
R90 a_2479_7336.n50 a_2479_7336.n37 8.28285
R91 a_2479_7336.n19 a_2479_7336.n6 8.28285
R92 a_2479_7336.n75 a_2479_7336.n64 8.22405
R93 a_2479_7336.n48 a_2479_7336.n36 6.77697
R94 a_2479_7336.n17 a_2479_7336.n5 6.77697
R95 a_2479_7336.n30 a_2479_7336.n28 6.19091
R96 a_2479_7336.n46 a_2479_7336.n35 5.27109
R97 a_2479_7336.n15 a_2479_7336.n4 5.27109
R98 a_2479_7336.n76 a_2479_7336.n75 4.66982
R99 a_2479_7336.n44 a_2479_7336.n34 3.76521
R100 a_2479_7336.n13 a_2479_7336.n3 3.76521
R101 a_2479_7336.n60 a_2479_7336.n59 3.31388
R102 a_2479_7336.n76 a_2479_7336.t14 2.8878
R103 a_2479_7336.n64 a_2479_7336.n62 2.87753
R104 a_2479_7336.n61 a_2479_7336.t13 2.48621
R105 a_2479_7336.n61 a_2479_7336.t5 2.48621
R106 a_2479_7336.n63 a_2479_7336.t4 2.48621
R107 a_2479_7336.n63 a_2479_7336.t2 2.48621
R108 a_2479_7336.n57 a_2479_7336.t6 2.48621
R109 a_2479_7336.n57 a_2479_7336.t8 2.48621
R110 a_2479_7336.n26 a_2479_7336.t11 2.48621
R111 a_2479_7336.n26 a_2479_7336.t3 2.48621
R112 a_2479_7336.n29 a_2479_7336.t15 2.48621
R113 a_2479_7336.n29 a_2479_7336.t12 2.48621
R114 a_2479_7336.n56 a_2479_7336.n55 2.36936
R115 a_2479_7336.n25 a_2479_7336.n24 2.36936
R116 a_2479_7336.n60 a_2479_7336.n30 2.30287
R117 a_2479_7336.n42 a_2479_7336.n33 2.25932
R118 a_2479_7336.n11 a_2479_7336.n2 2.25932
R119 a_2479_7336.n77 a_2479_7336.n76 1.41083
R120 a_2479_7336.n75 a_2479_7336.n74 1.3088
R121 a_2479_7336.n67 a_2479_7336.n66 0.3755
R122 a_2479_7336.n70 a_2479_7336.n69 0.3755
R123 a_2479_7336.n71 a_2479_7336.n70 0.3755
R124 a_2479_7336.n72 a_2479_7336.n71 0.3755
R125 a_2479_7336.n73 a_2479_7336.n72 0.3755
R126 a_2479_7336.n74 a_2479_7336.n73 0.3755
R127 a_2479_7336.n78 a_2479_7336.n77 0.3755
R128 a_2479_7336.n79 a_2479_7336.n78 0.3755
R129 a_2479_7336.n80 a_2479_7336.n79 0.3755
R130 a_2479_7336.n81 a_2479_7336.n80 0.3755
R131 a_2479_7336.n82 a_2479_7336.n81 0.3755
R132 a_2479_7336.n84 a_2479_7336.n83 0.3755
R133 a_2479_7336.n55 a_2479_7336.n41 0.320353
R134 a_2479_7336.n24 a_2479_7336.n10 0.320353
R135 a_2479_7336.n55 a_2479_7336.n54 0.196152
R136 a_2479_7336.n54 a_2479_7336.n53 0.196152
R137 a_2479_7336.n53 a_2479_7336.n51 0.196152
R138 a_2479_7336.n51 a_2479_7336.n49 0.196152
R139 a_2479_7336.n49 a_2479_7336.n47 0.196152
R140 a_2479_7336.n47 a_2479_7336.n45 0.196152
R141 a_2479_7336.n45 a_2479_7336.n43 0.196152
R142 a_2479_7336.n43 a_2479_7336.n31 0.196152
R143 a_2479_7336.n59 a_2479_7336.n31 0.196152
R144 a_2479_7336.n24 a_2479_7336.n23 0.196152
R145 a_2479_7336.n23 a_2479_7336.n22 0.196152
R146 a_2479_7336.n22 a_2479_7336.n20 0.196152
R147 a_2479_7336.n20 a_2479_7336.n18 0.196152
R148 a_2479_7336.n18 a_2479_7336.n16 0.196152
R149 a_2479_7336.n16 a_2479_7336.n14 0.196152
R150 a_2479_7336.n14 a_2479_7336.n12 0.196152
R151 a_2479_7336.n12 a_2479_7336.n0 0.196152
R152 a_2479_7336.n28 a_2479_7336.n0 0.196152
R153 a_2479_7336.n68 a_2479_7336.n67 0.188
R154 a_2479_7336.n69 a_2479_7336.n68 0.188
R155 a_2479_7336.n85 a_2479_7336.n82 0.188
R156 a_2479_7336.n85 a_2479_7336.n84 0.188
R157 VOUT.n31 VOUT.t26 260.298
R158 VOUT.t22 VOUT.n31 260.298
R159 VOUT.t26 VOUT.n26 260.298
R160 VOUT.n2 VOUT.t24 260.298
R161 VOUT.t20 VOUT.n2 260.298
R162 VOUT.n3 VOUT.t20 260.298
R163 VOUT.n32 VOUT.t22 260.111
R164 VOUT.t24 VOUT.n0 260.111
R165 VOUT.n30 VOUT.t28 232.03
R166 VOUT.t21 VOUT.n1 232.03
R167 VOUT.n20 VOUT.n18 206.708
R168 VOUT.n24 VOUT.n23 206.094
R169 VOUT.n22 VOUT.n21 206.094
R170 VOUT.n20 VOUT.n19 206.094
R171 VOUT.n16 VOUT.n15 206.094
R172 VOUT.n14 VOUT.n13 206.094
R173 VOUT.n12 VOUT.n11 206.094
R174 VOUT.n10 VOUT.n9 206.094
R175 VOUT.n29 VOUT.n28 203.03
R176 VOUT.n27 VOUT.n25 203.03
R177 VOUT.n7 VOUT.n6 203.03
R178 VOUT.n5 VOUT.n4 203.03
R179 VOUT.n62 VOUT.n61 185
R180 VOUT.n62 VOUT.n44 185
R181 VOUT.n62 VOUT.n43 185
R182 VOUT.n62 VOUT.n42 185
R183 VOUT.n62 VOUT.n41 185
R184 VOUT.n62 VOUT.n40 185
R185 VOUT.n62 VOUT.n39 185
R186 VOUT.n45 VOUT.t29 130.75
R187 VOUT.n45 VOUT.t31 91.3557
R188 VOUT.n63 VOUT.n62 86.5152
R189 VOUT.n47 VOUT.n38 30.3012
R190 VOUT.n28 VOUT.t23 28.5655
R191 VOUT.n28 VOUT.t27 28.5655
R192 VOUT.n27 VOUT.t14 28.5655
R193 VOUT.t23 VOUT.n27 28.5655
R194 VOUT.n23 VOUT.t3 28.5655
R195 VOUT.n23 VOUT.t16 28.5655
R196 VOUT.n21 VOUT.t7 28.5655
R197 VOUT.n21 VOUT.t12 28.5655
R198 VOUT.n19 VOUT.t2 28.5655
R199 VOUT.n19 VOUT.t15 28.5655
R200 VOUT.n18 VOUT.t10 28.5655
R201 VOUT.n18 VOUT.t11 28.5655
R202 VOUT.n6 VOUT.t25 28.5655
R203 VOUT.n6 VOUT.t8 28.5655
R204 VOUT.n5 VOUT.t21 28.5655
R205 VOUT.t25 VOUT.n5 28.5655
R206 VOUT.n15 VOUT.t13 28.5655
R207 VOUT.n15 VOUT.t1 28.5655
R208 VOUT.n13 VOUT.t0 28.5655
R209 VOUT.n13 VOUT.t5 28.5655
R210 VOUT.n11 VOUT.t17 28.5655
R211 VOUT.n11 VOUT.t6 28.5655
R212 VOUT.n9 VOUT.t9 28.5655
R213 VOUT.n9 VOUT.t4 28.5655
R214 VOUT.n61 VOUT.n37 24.8476
R215 VOUT.n60 VOUT.n44 23.3417
R216 VOUT.n64 VOUT.n63 22.0256
R217 VOUT.n57 VOUT.n43 21.8358
R218 VOUT.n55 VOUT.n42 20.3299
R219 VOUT.n65 VOUT.n64 19.0885
R220 VOUT.n53 VOUT.n41 18.824
R221 VOUT.n51 VOUT.n40 17.3181
R222 VOUT.n62 VOUT.n38 16.3559
R223 VOUT.n49 VOUT.n39 15.8123
R224 VOUT.n67 VOUT.t32 14.7991
R225 VOUT.n63 VOUT.n37 12.7256
R226 VOUT.n47 VOUT.n39 11.2946
R227 VOUT.n49 VOUT.n40 9.78874
R228 VOUT.n37 VOUT.n36 9.3005
R229 VOUT.n60 VOUT.n59 9.3005
R230 VOUT.n58 VOUT.n57 9.3005
R231 VOUT.n56 VOUT.n55 9.3005
R232 VOUT.n54 VOUT.n53 9.3005
R233 VOUT.n52 VOUT.n51 9.3005
R234 VOUT.n50 VOUT.n49 9.3005
R235 VOUT.n48 VOUT.n47 9.3005
R236 VOUT.n51 VOUT.n41 8.28285
R237 VOUT.n53 VOUT.n42 6.77697
R238 VOUT.n55 VOUT.n43 5.27109
R239 VOUT.t19 VOUT.n66 3.9533
R240 VOUT.n57 VOUT.n44 3.76521
R241 VOUT.n65 VOUT.n35 3.29996
R242 VOUT.n10 VOUT.n8 3.23261
R243 VOUT.n34 VOUT.n33 2.55612
R244 VOUT.n62 VOUT.t33 2.48621
R245 VOUT.n62 VOUT.t30 2.48621
R246 VOUT VOUT.n34 2.47337
R247 VOUT.n46 VOUT.n38 2.36936
R248 VOUT.n61 VOUT.n60 2.25932
R249 VOUT.n17 VOUT.n16 2.12962
R250 VOUT VOUT.n67 1.76033
R251 VOUT.n35 VOUT.n17 1.09816
R252 VOUT.n22 VOUT.n20 0.61449
R253 VOUT.n24 VOUT.n22 0.61449
R254 VOUT.n34 VOUT.n24 0.61449
R255 VOUT.n12 VOUT.n10 0.61449
R256 VOUT.n14 VOUT.n12 0.61449
R257 VOUT.n16 VOUT.n14 0.61449
R258 VOUT.n35 VOUT 0.521984
R259 VOUT.n8 VOUT.n7 0.446229
R260 VOUT.n7 VOUT.n1 0.43664
R261 VOUT.n30 VOUT.n25 0.436638
R262 VOUT.n33 VOUT.n25 0.38373
R263 VOUT.n29 VOUT.n26 0.38373
R264 VOUT.n4 VOUT.n3 0.383729
R265 VOUT.n46 VOUT.n45 0.320353
R266 VOUT.n31 VOUT.n30 0.285826
R267 VOUT.n2 VOUT.n1 0.285826
R268 VOUT.n66 VOUT.n65 0.220947
R269 VOUT.n64 VOUT.n36 0.196152
R270 VOUT.n59 VOUT.n36 0.196152
R271 VOUT.n59 VOUT.n58 0.196152
R272 VOUT.n58 VOUT.n56 0.196152
R273 VOUT.n56 VOUT.n54 0.196152
R274 VOUT.n54 VOUT.n52 0.196152
R275 VOUT.n52 VOUT.n50 0.196152
R276 VOUT.n50 VOUT.n48 0.196152
R277 VOUT.n48 VOUT.n46 0.196152
R278 VOUT.n33 VOUT.n32 0.188
R279 VOUT.n32 VOUT.n26 0.188
R280 VOUT.n3 VOUT.n0 0.188
R281 VOUT.n8 VOUT.n0 0.1255
R282 VOUT.n4 VOUT.n1 0.0984044
R283 VOUT.n30 VOUT.n29 0.0984028
R284 VOUT.n66 VOUT.n17 0.0649934
R285 VOUT.n67 VOUT.t19 0.0170587
R286 VOUT VOUT.t18 0.00167066
R287 VDD.n297 VDD.n68 723.529
R288 VDD.n73 VDD.n65 723.529
R289 VDD.n136 VDD.n112 723.529
R290 VDD.n180 VDD.n114 723.529
R291 VDD.n257 VDD.n256 515.294
R292 VDD.n55 VDD.n51 275.295
R293 VDD.n147 VDD.n131 275.295
R294 VDD.n34 VDD.t73 260.486
R295 VDD.n20 VDD.t52 260.486
R296 VDD.n330 VDD.t43 260.486
R297 VDD.n315 VDD.t58 260.486
R298 VDD.t38 VDD.n38 260.298
R299 VDD.n36 VDD.t54 260.298
R300 VDD.n39 VDD.t38 260.298
R301 VDD.t71 VDD.n19 260.298
R302 VDD.n17 VDD.t60 260.298
R303 VDD.n13 VDD.t60 260.298
R304 VDD.t47 VDD.n327 260.298
R305 VDD.t62 VDD.n329 260.298
R306 VDD.n334 VDD.t47 260.298
R307 VDD.n312 VDD.t69 260.298
R308 VDD.t69 VDD.n309 260.298
R309 VDD.n316 VDD.t75 260.298
R310 VDD.n1 VDD.t45 260.199
R311 VDD.n352 VDD.t64 260.199
R312 VDD.t56 VDD.n32 260.111
R313 VDD.n37 VDD.t56 260.111
R314 VDD.t54 VDD.n34 260.111
R315 VDD.n20 VDD.t71 260.111
R316 VDD.t41 VDD.n12 260.111
R317 VDD.n18 VDD.t41 260.111
R318 VDD.n333 VDD.t67 260.111
R319 VDD.t67 VDD.n332 260.111
R320 VDD.n330 VDD.t62 260.111
R321 VDD.t75 VDD.n315 260.111
R322 VDD.n314 VDD.t50 260.111
R323 VDD.t50 VDD.n313 260.111
R324 VDD.n67 VDD.n66 240
R325 VDD.n292 VDD.n66 240
R326 VDD.n290 VDD.n289 240
R327 VDD.n301 VDD.n50 240
R328 VDD.n253 VDD.n252 240
R329 VDD.n261 VDD.n260 240
R330 VDD.n265 VDD.n264 240
R331 VDD.n269 VDD.n268 240
R332 VDD.n273 VDD.n272 240
R333 VDD.n277 VDD.n276 240
R334 VDD.n279 VDD.n65 240
R335 VDD.n186 VDD.n112 240
R336 VDD.n186 VDD.n110 240
R337 VDD.n190 VDD.n110 240
R338 VDD.n190 VDD.n105 240
R339 VDD.n199 VDD.n105 240
R340 VDD.n199 VDD.n103 240
R341 VDD.n203 VDD.n103 240
R342 VDD.n203 VDD.n98 240
R343 VDD.n212 VDD.n98 240
R344 VDD.n212 VDD.n96 240
R345 VDD.n216 VDD.n96 240
R346 VDD.n216 VDD.n91 240
R347 VDD.n224 VDD.n91 240
R348 VDD.n224 VDD.n89 240
R349 VDD.n228 VDD.n89 240
R350 VDD.n228 VDD.n83 240
R351 VDD.n236 VDD.n83 240
R352 VDD.n236 VDD.n81 240
R353 VDD.n240 VDD.n81 240
R354 VDD.n240 VDD.n75 240
R355 VDD.n248 VDD.n75 240
R356 VDD.n248 VDD.n72 240
R357 VDD.n284 VDD.n72 240
R358 VDD.n284 VDD.n73 240
R359 VDD.n178 VDD.n177 240
R360 VDD.n175 VDD.n119 240
R361 VDD.n171 VDD.n170 240
R362 VDD.n168 VDD.n122 240
R363 VDD.n164 VDD.n163 240
R364 VDD.n161 VDD.n125 240
R365 VDD.n157 VDD.n156 240
R366 VDD.n154 VDD.n128 240
R367 VDD.n150 VDD.n149 240
R368 VDD.n143 VDD.n142 240
R369 VDD.n140 VDD.n134 240
R370 VDD.n184 VDD.n114 240
R371 VDD.n184 VDD.n109 240
R372 VDD.n193 VDD.n109 240
R373 VDD.n193 VDD.n107 240
R374 VDD.n197 VDD.n107 240
R375 VDD.n197 VDD.n102 240
R376 VDD.n206 VDD.n102 240
R377 VDD.n206 VDD.n100 240
R378 VDD.n210 VDD.n100 240
R379 VDD.n210 VDD.n95 240
R380 VDD.n218 VDD.n95 240
R381 VDD.n218 VDD.n93 240
R382 VDD.n222 VDD.n93 240
R383 VDD.n222 VDD.n87 240
R384 VDD.n230 VDD.n87 240
R385 VDD.n230 VDD.n85 240
R386 VDD.n234 VDD.n85 240
R387 VDD.n234 VDD.n79 240
R388 VDD.n242 VDD.n79 240
R389 VDD.n242 VDD.n77 240
R390 VDD.n246 VDD.n77 240
R391 VDD.n246 VDD.n70 240
R392 VDD.n286 VDD.n70 240
R393 VDD.n286 VDD.n68 240
R394 VDD.n31 VDD.t40 232.03
R395 VDD.n16 VDD.t61 232.03
R396 VDD.n335 VDD.t49 232.03
R397 VDD.t70 VDD.n308 232.03
R398 VDD.n351 VDD.t66 231.758
R399 VDD.n345 VDD.n343 206.48
R400 VDD.n324 VDD.n323 205.865
R401 VDD.n349 VDD.n348 205.865
R402 VDD.n347 VDD.n346 205.865
R403 VDD.n345 VDD.n344 205.865
R404 VDD.n9 VDD.n8 205.865
R405 VDD.n7 VDD.n6 205.865
R406 VDD.n5 VDD.n4 205.865
R407 VDD.n3 VDD.n2 205.865
R408 VDD.n28 VDD.n27 205.865
R409 VDD.n351 VDD.n350 203.143
R410 VDD.n45 VDD.n44 203.127
R411 VDD.n26 VDD.n25 203.127
R412 VDD.n341 VDD.n340 203.127
R413 VDD.n322 VDD.n321 203.127
R414 VDD.n43 VDD.n29 203.126
R415 VDD.n24 VDD.n10 203.126
R416 VDD.n339 VDD.n325 203.126
R417 VDD.n320 VDD.n306 203.126
R418 VDD.n42 VDD.n30 203.03
R419 VDD.n41 VDD.n40 203.03
R420 VDD.n23 VDD.n22 203.03
R421 VDD.n15 VDD.n14 203.03
R422 VDD.n338 VDD.n326 203.03
R423 VDD.n337 VDD.n336 203.03
R424 VDD.n319 VDD.n318 203.03
R425 VDD.n311 VDD.n310 203.03
R426 VDD.n182 VDD.n114 185
R427 VDD.n116 VDD.n114 185
R428 VDD.n184 VDD.n183 185
R429 VDD.n185 VDD.n184 185
R430 VDD.n109 VDD.n108 185
R431 VDD.n113 VDD.n109 185
R432 VDD.n194 VDD.n193 185
R433 VDD.n193 VDD.n192 185
R434 VDD.n195 VDD.n107 185
R435 VDD.n191 VDD.n107 185
R436 VDD.n197 VDD.n196 185
R437 VDD.n198 VDD.n197 185
R438 VDD.n102 VDD.n101 185
R439 VDD.n106 VDD.n102 185
R440 VDD.n207 VDD.n206 185
R441 VDD.n206 VDD.n205 185
R442 VDD.n208 VDD.n100 185
R443 VDD.n204 VDD.n100 185
R444 VDD.n210 VDD.n209 185
R445 VDD.n211 VDD.n210 185
R446 VDD.n95 VDD.n94 185
R447 VDD.n99 VDD.n95 185
R448 VDD.n219 VDD.n218 185
R449 VDD.n218 VDD.n217 185
R450 VDD.n220 VDD.n93 185
R451 VDD.n93 VDD.n92 185
R452 VDD.n222 VDD.n221 185
R453 VDD.n223 VDD.n222 185
R454 VDD.n87 VDD.n86 185
R455 VDD.n88 VDD.n87 185
R456 VDD.n231 VDD.n230 185
R457 VDD.n230 VDD.n229 185
R458 VDD.n232 VDD.n85 185
R459 VDD.n85 VDD.n84 185
R460 VDD.n234 VDD.n233 185
R461 VDD.n235 VDD.n234 185
R462 VDD.n79 VDD.n78 185
R463 VDD.n80 VDD.n79 185
R464 VDD.n243 VDD.n242 185
R465 VDD.n242 VDD.n241 185
R466 VDD.n244 VDD.n77 185
R467 VDD.n77 VDD.n76 185
R468 VDD.n246 VDD.n245 185
R469 VDD.n247 VDD.n246 185
R470 VDD.n70 VDD.n69 185
R471 VDD.n71 VDD.n70 185
R472 VDD.n287 VDD.n286 185
R473 VDD.n286 VDD.n285 185
R474 VDD.n288 VDD.n68 185
R475 VDD.n68 VDD.n52 185
R476 VDD.n137 VDD.n136 185
R477 VDD.n138 VDD.n134 185
R478 VDD.n140 VDD.n139 185
R479 VDD.n142 VDD.n132 185
R480 VDD.n144 VDD.n143 185
R481 VDD.n145 VDD.n131 185
R482 VDD.n147 VDD.n146 185
R483 VDD.n149 VDD.n129 185
R484 VDD.n151 VDD.n150 185
R485 VDD.n152 VDD.n128 185
R486 VDD.n154 VDD.n153 185
R487 VDD.n156 VDD.n126 185
R488 VDD.n158 VDD.n157 185
R489 VDD.n159 VDD.n125 185
R490 VDD.n161 VDD.n160 185
R491 VDD.n163 VDD.n123 185
R492 VDD.n165 VDD.n164 185
R493 VDD.n166 VDD.n122 185
R494 VDD.n168 VDD.n167 185
R495 VDD.n170 VDD.n120 185
R496 VDD.n172 VDD.n171 185
R497 VDD.n173 VDD.n119 185
R498 VDD.n175 VDD.n174 185
R499 VDD.n177 VDD.n118 185
R500 VDD.n178 VDD.n115 185
R501 VDD.n181 VDD.n180 185
R502 VDD.n282 VDD.n73 185
R503 VDD.n73 VDD.n52 185
R504 VDD.n284 VDD.n283 185
R505 VDD.n285 VDD.n284 185
R506 VDD.n250 VDD.n72 185
R507 VDD.n72 VDD.n71 185
R508 VDD.n249 VDD.n248 185
R509 VDD.n248 VDD.n247 185
R510 VDD.n75 VDD.n74 185
R511 VDD.n76 VDD.n75 185
R512 VDD.n240 VDD.n239 185
R513 VDD.n241 VDD.n240 185
R514 VDD.n238 VDD.n81 185
R515 VDD.n81 VDD.n80 185
R516 VDD.n237 VDD.n236 185
R517 VDD.n236 VDD.n235 185
R518 VDD.n83 VDD.n82 185
R519 VDD.n84 VDD.n83 185
R520 VDD.n228 VDD.n227 185
R521 VDD.n229 VDD.n228 185
R522 VDD.n226 VDD.n89 185
R523 VDD.n89 VDD.n88 185
R524 VDD.n225 VDD.n224 185
R525 VDD.n224 VDD.n223 185
R526 VDD.n91 VDD.n90 185
R527 VDD.n92 VDD.n91 185
R528 VDD.n216 VDD.n215 185
R529 VDD.n217 VDD.n216 185
R530 VDD.n214 VDD.n96 185
R531 VDD.n99 VDD.n96 185
R532 VDD.n213 VDD.n212 185
R533 VDD.n212 VDD.n211 185
R534 VDD.n98 VDD.n97 185
R535 VDD.n204 VDD.n98 185
R536 VDD.n203 VDD.n202 185
R537 VDD.n205 VDD.n203 185
R538 VDD.n201 VDD.n103 185
R539 VDD.n106 VDD.n103 185
R540 VDD.n200 VDD.n199 185
R541 VDD.n199 VDD.n198 185
R542 VDD.n105 VDD.n104 185
R543 VDD.n191 VDD.n105 185
R544 VDD.n190 VDD.n189 185
R545 VDD.n192 VDD.n190 185
R546 VDD.n188 VDD.n110 185
R547 VDD.n113 VDD.n110 185
R548 VDD.n187 VDD.n186 185
R549 VDD.n186 VDD.n185 185
R550 VDD.n112 VDD.n111 185
R551 VDD.n116 VDD.n112 185
R552 VDD.n297 VDD.n296 185
R553 VDD.n295 VDD.n67 185
R554 VDD.n294 VDD.n66 185
R555 VDD.n299 VDD.n66 185
R556 VDD.n293 VDD.n292 185
R557 VDD.n291 VDD.n290 185
R558 VDD.n289 VDD.n47 185
R559 VDD.n55 VDD.n54 185
R560 VDD.n51 VDD.n48 185
R561 VDD.n302 VDD.n301 185
R562 VDD.n50 VDD.n49 185
R563 VDD.n252 VDD.n251 185
R564 VDD.n254 VDD.n253 185
R565 VDD.n256 VDD.n255 185
R566 VDD.n258 VDD.n257 185
R567 VDD.n260 VDD.n259 185
R568 VDD.n262 VDD.n261 185
R569 VDD.n264 VDD.n263 185
R570 VDD.n266 VDD.n265 185
R571 VDD.n268 VDD.n267 185
R572 VDD.n270 VDD.n269 185
R573 VDD.n272 VDD.n271 185
R574 VDD.n274 VDD.n273 185
R575 VDD.n276 VDD.n275 185
R576 VDD.n278 VDD.n277 185
R577 VDD.n280 VDD.n279 185
R578 VDD.n281 VDD.n65 185
R579 VDD.n299 VDD.n65 185
R580 VDD.n157 VDD.n127 107.683
R581 VDD.n127 VDD.n125 107.683
R582 VDD.n1 VDD.n0 101.662
R583 VDD.n269 VDD.n62 78.9253
R584 VDD.n169 VDD.n168 78.9253
R585 VDD.n170 VDD.n169 78.9253
R586 VDD.n272 VDD.n62 78.9253
R587 VDD.n182 VDD.n181 77.177
R588 VDD.n296 VDD.n288 77.177
R589 VDD.n137 VDD.n111 77.177
R590 VDD.n282 VDD.n281 77.177
R591 VDD.n298 VDD.n297 72.7879
R592 VDD.n292 VDD.n53 72.7879
R593 VDD.n289 VDD.n56 72.7879
R594 VDD.n300 VDD.n51 72.7879
R595 VDD.n57 VDD.n50 72.7879
R596 VDD.n253 VDD.n58 72.7879
R597 VDD.n257 VDD.n59 72.7879
R598 VDD.n261 VDD.n60 72.7879
R599 VDD.n265 VDD.n61 72.7879
R600 VDD.n273 VDD.n63 72.7879
R601 VDD.n277 VDD.n64 72.7879
R602 VDD.n179 VDD.n178 72.7879
R603 VDD.n176 VDD.n175 72.7879
R604 VDD.n171 VDD.n121 72.7879
R605 VDD.n164 VDD.n124 72.7879
R606 VDD.n162 VDD.n161 72.7879
R607 VDD.n155 VDD.n154 72.7879
R608 VDD.n150 VDD.n130 72.7879
R609 VDD.n148 VDD.n147 72.7879
R610 VDD.n143 VDD.n133 72.7879
R611 VDD.n141 VDD.n140 72.7879
R612 VDD.n136 VDD.n135 72.7879
R613 VDD.n135 VDD.n134 72.7879
R614 VDD.n142 VDD.n141 72.7879
R615 VDD.n133 VDD.n131 72.7879
R616 VDD.n149 VDD.n148 72.7879
R617 VDD.n130 VDD.n128 72.7879
R618 VDD.n156 VDD.n155 72.7879
R619 VDD.n163 VDD.n162 72.7879
R620 VDD.n124 VDD.n122 72.7879
R621 VDD.n121 VDD.n119 72.7879
R622 VDD.n177 VDD.n176 72.7879
R623 VDD.n180 VDD.n179 72.7879
R624 VDD.n298 VDD.n67 72.7879
R625 VDD.n290 VDD.n53 72.7879
R626 VDD.n56 VDD.n55 72.7879
R627 VDD.n301 VDD.n300 72.7879
R628 VDD.n252 VDD.n57 72.7879
R629 VDD.n256 VDD.n58 72.7879
R630 VDD.n260 VDD.n59 72.7879
R631 VDD.n264 VDD.n60 72.7879
R632 VDD.n268 VDD.n61 72.7879
R633 VDD.n276 VDD.n63 72.7879
R634 VDD.n279 VDD.n64 72.7879
R635 VDD.n117 VDD.n116 57.1093
R636 VDD.n299 VDD.n52 57.1093
R637 VDD.n135 VDD.n117 56.1076
R638 VDD.n141 VDD.n117 56.1076
R639 VDD.n133 VDD.n117 56.1076
R640 VDD.n148 VDD.n117 56.1076
R641 VDD.n130 VDD.n117 56.1076
R642 VDD.n155 VDD.n117 56.1076
R643 VDD.n162 VDD.n117 56.1076
R644 VDD.n124 VDD.n117 56.1076
R645 VDD.n121 VDD.n117 56.1076
R646 VDD.n176 VDD.n117 56.1076
R647 VDD.n179 VDD.n117 56.1076
R648 VDD.n299 VDD.n298 56.1076
R649 VDD.n299 VDD.n53 56.1076
R650 VDD.n299 VDD.n56 56.1076
R651 VDD.n300 VDD.n299 56.1076
R652 VDD.n299 VDD.n57 56.1076
R653 VDD.n299 VDD.n58 56.1076
R654 VDD.n299 VDD.n59 56.1076
R655 VDD.n299 VDD.n60 56.1076
R656 VDD.n299 VDD.n61 56.1076
R657 VDD.n299 VDD.n63 56.1076
R658 VDD.n299 VDD.n64 56.1076
R659 VDD.n159 VDD.n158 54.9652
R660 VDD.n258 VDD.n255 54.9652
R661 VDD.n169 VDD.n117 53.0388
R662 VDD.n299 VDD.n62 53.0388
R663 VDD.n0 VDD.t22 41.0864
R664 VDD.n127 VDD.n117 38.6605
R665 VDD.n185 VDD.n113 30.8211
R666 VDD.n192 VDD.n191 30.8211
R667 VDD.n198 VDD.n106 30.8211
R668 VDD.n205 VDD.n204 30.8211
R669 VDD.n211 VDD.n99 30.8211
R670 VDD.n217 VDD.n92 30.8211
R671 VDD.n223 VDD.n92 30.8211
R672 VDD.n229 VDD.n88 30.8211
R673 VDD.n235 VDD.n84 30.8211
R674 VDD.n241 VDD.n80 30.8211
R675 VDD.n247 VDD.n76 30.8211
R676 VDD.n285 VDD.n71 30.8211
R677 VDD.n99 VDD.t18 30.3679
R678 VDD.t2 VDD.n88 30.3679
R679 VDD.n204 VDD.t5 29.4614
R680 VDD.t0 VDD.n84 29.4614
R681 VDD.n167 VDD.n120 29.3652
R682 VDD.n146 VDD.n145 29.3652
R683 VDD.n54 VDD.n48 29.3652
R684 VDD.n271 VDD.n270 29.3652
R685 VDD.n8 VDD.t17 28.5655
R686 VDD.n8 VDD.t30 28.5655
R687 VDD.n6 VDD.t11 28.5655
R688 VDD.n6 VDD.t7 28.5655
R689 VDD.n4 VDD.t24 28.5655
R690 VDD.n4 VDD.t20 28.5655
R691 VDD.n2 VDD.t14 28.5655
R692 VDD.n2 VDD.t29 28.5655
R693 VDD.t55 VDD.n42 28.5655
R694 VDD.n42 VDD.t57 28.5655
R695 VDD.t57 VDD.n41 28.5655
R696 VDD.n41 VDD.t39 28.5655
R697 VDD.t74 VDD.n43 28.5655
R698 VDD.n43 VDD.t55 28.5655
R699 VDD.n44 VDD.t1 28.5655
R700 VDD.n44 VDD.t74 28.5655
R701 VDD.n27 VDD.t36 28.5655
R702 VDD.n27 VDD.t3 28.5655
R703 VDD.n23 VDD.t42 28.5655
R704 VDD.t72 VDD.n23 28.5655
R705 VDD.n14 VDD.t61 28.5655
R706 VDD.n14 VDD.t42 28.5655
R707 VDD.n24 VDD.t72 28.5655
R708 VDD.t53 VDD.n24 28.5655
R709 VDD.n25 VDD.t53 28.5655
R710 VDD.n25 VDD.t6 28.5655
R711 VDD.n340 VDD.t4 28.5655
R712 VDD.n340 VDD.t44 28.5655
R713 VDD.t63 VDD.n338 28.5655
R714 VDD.n338 VDD.t68 28.5655
R715 VDD.t68 VDD.n337 28.5655
R716 VDD.n337 VDD.t48 28.5655
R717 VDD.t44 VDD.n339 28.5655
R718 VDD.n339 VDD.t63 28.5655
R719 VDD.n321 VDD.t59 28.5655
R720 VDD.n321 VDD.t37 28.5655
R721 VDD.n319 VDD.t51 28.5655
R722 VDD.t76 VDD.n319 28.5655
R723 VDD.n310 VDD.t70 28.5655
R724 VDD.n310 VDD.t51 28.5655
R725 VDD.n320 VDD.t76 28.5655
R726 VDD.t59 VDD.n320 28.5655
R727 VDD.n323 VDD.t35 28.5655
R728 VDD.n323 VDD.t34 28.5655
R729 VDD.n350 VDD.t9 28.5655
R730 VDD.n350 VDD.t65 28.5655
R731 VDD.n348 VDD.t16 28.5655
R732 VDD.n348 VDD.t28 28.5655
R733 VDD.n346 VDD.t10 28.5655
R734 VDD.n346 VDD.t31 28.5655
R735 VDD.n344 VDD.t23 28.5655
R736 VDD.n344 VDD.t19 28.5655
R737 VDD.n343 VDD.t13 28.5655
R738 VDD.n343 VDD.t26 28.5655
R739 VDD.n106 VDD.t25 28.5549
R740 VDD.t15 VDD.n80 28.5549
R741 VDD.n191 VDD.t12 27.6484
R742 VDD.t27 VDD.n76 27.6484
R743 VDD.n113 VDD.t21 26.7419
R744 VDD.t8 VDD.n71 26.7419
R745 VDD.n116 VDD.t32 25.8354
R746 VDD.t33 VDD.n52 25.8354
R747 VDD.n183 VDD.n182 25.6005
R748 VDD.n183 VDD.n108 25.6005
R749 VDD.n194 VDD.n108 25.6005
R750 VDD.n195 VDD.n194 25.6005
R751 VDD.n196 VDD.n195 25.6005
R752 VDD.n196 VDD.n101 25.6005
R753 VDD.n207 VDD.n101 25.6005
R754 VDD.n208 VDD.n207 25.6005
R755 VDD.n209 VDD.n208 25.6005
R756 VDD.n209 VDD.n94 25.6005
R757 VDD.n219 VDD.n94 25.6005
R758 VDD.n220 VDD.n219 25.6005
R759 VDD.n221 VDD.n220 25.6005
R760 VDD.n221 VDD.n86 25.6005
R761 VDD.n231 VDD.n86 25.6005
R762 VDD.n232 VDD.n231 25.6005
R763 VDD.n233 VDD.n232 25.6005
R764 VDD.n233 VDD.n78 25.6005
R765 VDD.n243 VDD.n78 25.6005
R766 VDD.n244 VDD.n243 25.6005
R767 VDD.n245 VDD.n244 25.6005
R768 VDD.n245 VDD.n69 25.6005
R769 VDD.n287 VDD.n69 25.6005
R770 VDD.n288 VDD.n287 25.6005
R771 VDD.n181 VDD.n115 25.6005
R772 VDD.n118 VDD.n115 25.6005
R773 VDD.n174 VDD.n118 25.6005
R774 VDD.n174 VDD.n173 25.6005
R775 VDD.n173 VDD.n172 25.6005
R776 VDD.n172 VDD.n120 25.6005
R777 VDD.n167 VDD.n166 25.6005
R778 VDD.n166 VDD.n165 25.6005
R779 VDD.n165 VDD.n123 25.6005
R780 VDD.n160 VDD.n123 25.6005
R781 VDD.n160 VDD.n159 25.6005
R782 VDD.n158 VDD.n126 25.6005
R783 VDD.n153 VDD.n126 25.6005
R784 VDD.n153 VDD.n152 25.6005
R785 VDD.n152 VDD.n151 25.6005
R786 VDD.n151 VDD.n129 25.6005
R787 VDD.n146 VDD.n129 25.6005
R788 VDD.n145 VDD.n144 25.6005
R789 VDD.n144 VDD.n132 25.6005
R790 VDD.n139 VDD.n132 25.6005
R791 VDD.n139 VDD.n138 25.6005
R792 VDD.n138 VDD.n137 25.6005
R793 VDD.n187 VDD.n111 25.6005
R794 VDD.n188 VDD.n187 25.6005
R795 VDD.n189 VDD.n188 25.6005
R796 VDD.n189 VDD.n104 25.6005
R797 VDD.n200 VDD.n104 25.6005
R798 VDD.n201 VDD.n200 25.6005
R799 VDD.n202 VDD.n201 25.6005
R800 VDD.n202 VDD.n97 25.6005
R801 VDD.n213 VDD.n97 25.6005
R802 VDD.n214 VDD.n213 25.6005
R803 VDD.n215 VDD.n214 25.6005
R804 VDD.n215 VDD.n90 25.6005
R805 VDD.n225 VDD.n90 25.6005
R806 VDD.n226 VDD.n225 25.6005
R807 VDD.n227 VDD.n226 25.6005
R808 VDD.n227 VDD.n82 25.6005
R809 VDD.n237 VDD.n82 25.6005
R810 VDD.n238 VDD.n237 25.6005
R811 VDD.n239 VDD.n238 25.6005
R812 VDD.n239 VDD.n74 25.6005
R813 VDD.n249 VDD.n74 25.6005
R814 VDD.n250 VDD.n249 25.6005
R815 VDD.n283 VDD.n250 25.6005
R816 VDD.n283 VDD.n282 25.6005
R817 VDD.n296 VDD.n295 25.6005
R818 VDD.n295 VDD.n294 25.6005
R819 VDD.n294 VDD.n293 25.6005
R820 VDD.n293 VDD.n291 25.6005
R821 VDD.n291 VDD.n47 25.6005
R822 VDD.n54 VDD.n47 25.6005
R823 VDD.n302 VDD.n49 25.6005
R824 VDD.n251 VDD.n49 25.6005
R825 VDD.n254 VDD.n251 25.6005
R826 VDD.n255 VDD.n254 25.6005
R827 VDD.n259 VDD.n258 25.6005
R828 VDD.n262 VDD.n259 25.6005
R829 VDD.n263 VDD.n262 25.6005
R830 VDD.n266 VDD.n263 25.6005
R831 VDD.n267 VDD.n266 25.6005
R832 VDD.n270 VDD.n267 25.6005
R833 VDD.n274 VDD.n271 25.6005
R834 VDD.n275 VDD.n274 25.6005
R835 VDD.n278 VDD.n275 25.6005
R836 VDD.n280 VDD.n278 25.6005
R837 VDD.n281 VDD.n280 25.6005
R838 VDD.n303 VDD.n302 23.3417
R839 VDD.n0 VDD.t46 14.285
R840 VDD.n304 VDD.n303 9.3686
R841 VDD.n304 VDD.n47 9.36343
R842 VDD.n185 VDD.t32 4.98619
R843 VDD.n285 VDD.t33 4.98619
R844 VDD.n192 VDD.t21 4.0797
R845 VDD.n247 VDD.t8 4.0797
R846 VDD.n28 VDD.n26 3.35217
R847 VDD.n324 VDD.n322 3.35217
R848 VDD.n198 VDD.t12 3.17321
R849 VDD.n241 VDD.t27 3.17321
R850 VDD.n3 VDD.n1 3.06997
R851 VDD.n46 VDD.n45 2.73818
R852 VDD.n342 VDD.n341 2.73818
R853 VDD VDD.n356 2.72726
R854 VDD.n353 VDD.n352 2.45598
R855 VDD.n205 VDD.t25 2.26672
R856 VDD.n235 VDD.t15 2.26672
R857 VDD.n303 VDD.n48 2.25932
R858 VDD.n305 VDD.n304 2.20937
R859 VDD.n354 VDD.n342 2.07758
R860 VDD.n356 VDD.n9 1.76955
R861 VDD.n354 VDD.n353 1.63948
R862 VDD.n305 VDD.n46 1.485
R863 VDD.n211 VDD.t5 1.36023
R864 VDD.n229 VDD.t0 1.36023
R865 VDD.n355 VDD.n354 0.9725
R866 VDD.n5 VDD.n3 0.61449
R867 VDD.n7 VDD.n5 0.61449
R868 VDD.n9 VDD.n7 0.61449
R869 VDD.n46 VDD.n28 0.61449
R870 VDD.n342 VDD.n324 0.61449
R871 VDD.n347 VDD.n345 0.61449
R872 VDD.n349 VDD.n347 0.61449
R873 VDD.n353 VDD.n349 0.61449
R874 VDD.n355 VDD.n305 0.590949
R875 VDD.n356 VDD.n355 0.4865
R876 VDD.n217 VDD.t18 0.453744
R877 VDD.n223 VDD.t2 0.453744
R878 VDD.n336 VDD.n327 0.38373
R879 VDD.n331 VDD.n326 0.38373
R880 VDD.n312 VDD.n311 0.38373
R881 VDD.n318 VDD.n307 0.38373
R882 VDD.n40 VDD.n39 0.383729
R883 VDD.n33 VDD.n30 0.383729
R884 VDD.n15 VDD.n13 0.383729
R885 VDD.n22 VDD.n21 0.383729
R886 VDD.n35 VDD.n31 0.338735
R887 VDD.n35 VDD.n29 0.338735
R888 VDD.n45 VDD.n29 0.338735
R889 VDD.n16 VDD.n11 0.338735
R890 VDD.n11 VDD.n10 0.338735
R891 VDD.n26 VDD.n10 0.338735
R892 VDD.n335 VDD.n328 0.338735
R893 VDD.n328 VDD.n325 0.338735
R894 VDD.n341 VDD.n325 0.338735
R895 VDD.n317 VDD.n308 0.338735
R896 VDD.n317 VDD.n306 0.338735
R897 VDD.n322 VDD.n306 0.338735
R898 VDD.n38 VDD.n31 0.285826
R899 VDD.n36 VDD.n35 0.285826
R900 VDD.n17 VDD.n16 0.285826
R901 VDD.n19 VDD.n11 0.285826
R902 VDD.n335 VDD.n334 0.285826
R903 VDD.n329 VDD.n328 0.285826
R904 VDD.n309 VDD.n308 0.285826
R905 VDD.n317 VDD.n316 0.285826
R906 VDD.n37 VDD.n36 0.188
R907 VDD.n38 VDD.n37 0.188
R908 VDD.n34 VDD.n33 0.188
R909 VDD.n33 VDD.n32 0.188
R910 VDD.n39 VDD.n32 0.188
R911 VDD.n18 VDD.n17 0.188
R912 VDD.n19 VDD.n18 0.188
R913 VDD.n13 VDD.n12 0.188
R914 VDD.n21 VDD.n12 0.188
R915 VDD.n21 VDD.n20 0.188
R916 VDD.n331 VDD.n330 0.188
R917 VDD.n332 VDD.n331 0.188
R918 VDD.n332 VDD.n327 0.188
R919 VDD.n333 VDD.n329 0.188
R920 VDD.n334 VDD.n333 0.188
R921 VDD.n313 VDD.n312 0.188
R922 VDD.n313 VDD.n307 0.188
R923 VDD.n315 VDD.n307 0.188
R924 VDD.n314 VDD.n309 0.188
R925 VDD.n316 VDD.n314 0.188
R926 VDD.n40 VDD.n31 0.0984044
R927 VDD.n35 VDD.n30 0.0984044
R928 VDD.n16 VDD.n15 0.0984044
R929 VDD.n22 VDD.n11 0.0984044
R930 VDD.n328 VDD.n326 0.0984028
R931 VDD.n336 VDD.n335 0.0984028
R932 VDD.n318 VDD.n317 0.0984028
R933 VDD.n311 VDD.n308 0.0984028
R934 VDD.n352 VDD.n351 0.0793043
R935 VSS.n1463 VSS.n617 5684.63
R936 VSS.n2117 VSS.n642 1321.06
R937 VSS.n2119 VSS.n640 1321.06
R938 VSS.n2286 VSS.n530 1321.06
R939 VSS.n2278 VSS.n2277 1321.06
R940 VSS.n1786 VSS.n856 1268.91
R941 VSS.n1867 VSS.n836 1268.91
R942 VSS.n1742 VSS.n1741 1268.91
R943 VSS.n1820 VSS.n834 1268.91
R944 VSS.n1293 VSS.n1236 1268.91
R945 VSS.n1589 VSS.n1093 1268.91
R946 VSS.n1295 VSS.n1235 1268.91
R947 VSS.n1546 VSS.n1545 1268.91
R948 VSS.n1608 VSS.n1023 1268.91
R949 VSS.n1715 VSS.n881 1268.91
R950 VSS.n1672 VSS.n1671 1268.91
R951 VSS.n1610 VSS.n1020 1268.91
R952 VSS.n516 VSS.n260 1182
R953 VSS.n2540 VSS.n142 1182
R954 VSS.n514 VSS.n262 1182
R955 VSS.n2484 VSS.n147 1182
R956 VSS.n1466 VSS.n1119 1182
R957 VSS.n2067 VSS.n768 1182
R958 VSS.n1331 VSS.n1330 1182
R959 VSS.n1880 VSS.n818 1182
R960 VSS.n2023 VSS.n822 996.588
R961 VSS.n1975 VSS.n1974 602.588
R962 VSS.n1927 VSS.n1926 602.588
R963 VSS.n2120 VSS.n2119 585
R964 VSS.n2119 VSS.n2118 585
R965 VSS.n2121 VSS.n638 585
R966 VSS.n638 VSS.n637 585
R967 VSS.n2123 VSS.n2122 585
R968 VSS.n2124 VSS.n2123 585
R969 VSS.n632 VSS.n631 585
R970 VSS.n633 VSS.n632 585
R971 VSS.n2132 VSS.n2131 585
R972 VSS.n2131 VSS.n2130 585
R973 VSS.n2133 VSS.n630 585
R974 VSS.n630 VSS.n629 585
R975 VSS.n2135 VSS.n2134 585
R976 VSS.n2136 VSS.n2135 585
R977 VSS.n624 VSS.n623 585
R978 VSS.n625 VSS.n624 585
R979 VSS.n2144 VSS.n2143 585
R980 VSS.n2143 VSS.n2142 585
R981 VSS.n2145 VSS.n622 585
R982 VSS.n622 VSS.n621 585
R983 VSS.n2147 VSS.n2146 585
R984 VSS.n2148 VSS.n2147 585
R985 VSS.n615 VSS.n614 585
R986 VSS.n616 VSS.n615 585
R987 VSS.n2156 VSS.n2155 585
R988 VSS.n2155 VSS.n2154 585
R989 VSS.n2157 VSS.n613 585
R990 VSS.n613 VSS.n612 585
R991 VSS.n2159 VSS.n2158 585
R992 VSS.n2160 VSS.n2159 585
R993 VSS.n607 VSS.n606 585
R994 VSS.n608 VSS.n607 585
R995 VSS.n2168 VSS.n2167 585
R996 VSS.n2167 VSS.n2166 585
R997 VSS.n2169 VSS.n605 585
R998 VSS.n605 VSS.n604 585
R999 VSS.n2171 VSS.n2170 585
R1000 VSS.n2172 VSS.n2171 585
R1001 VSS.n599 VSS.n598 585
R1002 VSS.n600 VSS.n599 585
R1003 VSS.n2180 VSS.n2179 585
R1004 VSS.n2179 VSS.n2178 585
R1005 VSS.n2181 VSS.n597 585
R1006 VSS.n597 VSS.n596 585
R1007 VSS.n2183 VSS.n2182 585
R1008 VSS.n2184 VSS.n2183 585
R1009 VSS.n591 VSS.n590 585
R1010 VSS.n592 VSS.n591 585
R1011 VSS.n2192 VSS.n2191 585
R1012 VSS.n2191 VSS.n2190 585
R1013 VSS.n2193 VSS.n589 585
R1014 VSS.n589 VSS.n588 585
R1015 VSS.n2195 VSS.n2194 585
R1016 VSS.n2196 VSS.n2195 585
R1017 VSS.n583 VSS.n582 585
R1018 VSS.n584 VSS.n583 585
R1019 VSS.n2204 VSS.n2203 585
R1020 VSS.n2203 VSS.n2202 585
R1021 VSS.n2205 VSS.n581 585
R1022 VSS.n581 VSS.n580 585
R1023 VSS.n2207 VSS.n2206 585
R1024 VSS.n2208 VSS.n2207 585
R1025 VSS.n575 VSS.n574 585
R1026 VSS.n576 VSS.n575 585
R1027 VSS.n2216 VSS.n2215 585
R1028 VSS.n2215 VSS.n2214 585
R1029 VSS.n2217 VSS.n573 585
R1030 VSS.n573 VSS.n572 585
R1031 VSS.n2219 VSS.n2218 585
R1032 VSS.n2220 VSS.n2219 585
R1033 VSS.n567 VSS.n566 585
R1034 VSS.n568 VSS.n567 585
R1035 VSS.n2228 VSS.n2227 585
R1036 VSS.n2227 VSS.n2226 585
R1037 VSS.n2229 VSS.n565 585
R1038 VSS.n565 VSS.n564 585
R1039 VSS.n2231 VSS.n2230 585
R1040 VSS.n2232 VSS.n2231 585
R1041 VSS.n559 VSS.n558 585
R1042 VSS.n560 VSS.n559 585
R1043 VSS.n2240 VSS.n2239 585
R1044 VSS.n2239 VSS.n2238 585
R1045 VSS.n2241 VSS.n557 585
R1046 VSS.n557 VSS.n556 585
R1047 VSS.n2243 VSS.n2242 585
R1048 VSS.n2244 VSS.n2243 585
R1049 VSS.n551 VSS.n550 585
R1050 VSS.n552 VSS.n551 585
R1051 VSS.n2252 VSS.n2251 585
R1052 VSS.n2251 VSS.n2250 585
R1053 VSS.n2253 VSS.n549 585
R1054 VSS.n549 VSS.n548 585
R1055 VSS.n2255 VSS.n2254 585
R1056 VSS.n2256 VSS.n2255 585
R1057 VSS.n543 VSS.n542 585
R1058 VSS.n544 VSS.n543 585
R1059 VSS.n2264 VSS.n2263 585
R1060 VSS.n2263 VSS.n2262 585
R1061 VSS.n2265 VSS.n541 585
R1062 VSS.n541 VSS.n540 585
R1063 VSS.n2268 VSS.n2267 585
R1064 VSS.n2269 VSS.n2268 585
R1065 VSS.n2266 VSS.n534 585
R1066 VSS.n536 VSS.n534 585
R1067 VSS.n2276 VSS.n535 585
R1068 VSS.n2276 VSS.n2275 585
R1069 VSS.n2277 VSS.n533 585
R1070 VSS.n2277 VSS.n527 585
R1071 VSS.n2279 VSS.n2278 585
R1072 VSS.n2281 VSS.n2280 585
R1073 VSS.n2283 VSS.n2282 585
R1074 VSS.n2284 VSS.n531 585
R1075 VSS.n2286 VSS.n2285 585
R1076 VSS.n2287 VSS.n2286 585
R1077 VSS.n532 VSS.n530 585
R1078 VSS.n530 VSS.n527 585
R1079 VSS.n2274 VSS.n2273 585
R1080 VSS.n2275 VSS.n2274 585
R1081 VSS.n2272 VSS.n537 585
R1082 VSS.n537 VSS.n536 585
R1083 VSS.n2271 VSS.n2270 585
R1084 VSS.n2270 VSS.n2269 585
R1085 VSS.n539 VSS.n538 585
R1086 VSS.n540 VSS.n539 585
R1087 VSS.n2261 VSS.n2260 585
R1088 VSS.n2262 VSS.n2261 585
R1089 VSS.n2259 VSS.n545 585
R1090 VSS.n545 VSS.n544 585
R1091 VSS.n2258 VSS.n2257 585
R1092 VSS.n2257 VSS.n2256 585
R1093 VSS.n547 VSS.n546 585
R1094 VSS.n548 VSS.n547 585
R1095 VSS.n2249 VSS.n2248 585
R1096 VSS.n2250 VSS.n2249 585
R1097 VSS.n2247 VSS.n553 585
R1098 VSS.n553 VSS.n552 585
R1099 VSS.n2246 VSS.n2245 585
R1100 VSS.n2245 VSS.n2244 585
R1101 VSS.n555 VSS.n554 585
R1102 VSS.n556 VSS.n555 585
R1103 VSS.n2237 VSS.n2236 585
R1104 VSS.n2238 VSS.n2237 585
R1105 VSS.n2235 VSS.n561 585
R1106 VSS.n561 VSS.n560 585
R1107 VSS.n2234 VSS.n2233 585
R1108 VSS.n2233 VSS.n2232 585
R1109 VSS.n563 VSS.n562 585
R1110 VSS.n564 VSS.n563 585
R1111 VSS.n2225 VSS.n2224 585
R1112 VSS.n2226 VSS.n2225 585
R1113 VSS.n2223 VSS.n569 585
R1114 VSS.n569 VSS.n568 585
R1115 VSS.n2222 VSS.n2221 585
R1116 VSS.n2221 VSS.n2220 585
R1117 VSS.n571 VSS.n570 585
R1118 VSS.n572 VSS.n571 585
R1119 VSS.n2213 VSS.n2212 585
R1120 VSS.n2214 VSS.n2213 585
R1121 VSS.n2211 VSS.n577 585
R1122 VSS.n577 VSS.n576 585
R1123 VSS.n2210 VSS.n2209 585
R1124 VSS.n2209 VSS.n2208 585
R1125 VSS.n579 VSS.n578 585
R1126 VSS.n580 VSS.n579 585
R1127 VSS.n2201 VSS.n2200 585
R1128 VSS.n2202 VSS.n2201 585
R1129 VSS.n2199 VSS.n585 585
R1130 VSS.n585 VSS.n584 585
R1131 VSS.n2198 VSS.n2197 585
R1132 VSS.n2197 VSS.n2196 585
R1133 VSS.n587 VSS.n586 585
R1134 VSS.n588 VSS.n587 585
R1135 VSS.n2189 VSS.n2188 585
R1136 VSS.n2190 VSS.n2189 585
R1137 VSS.n2187 VSS.n593 585
R1138 VSS.n593 VSS.n592 585
R1139 VSS.n2186 VSS.n2185 585
R1140 VSS.n2185 VSS.n2184 585
R1141 VSS.n595 VSS.n594 585
R1142 VSS.n596 VSS.n595 585
R1143 VSS.n2177 VSS.n2176 585
R1144 VSS.n2178 VSS.n2177 585
R1145 VSS.n2175 VSS.n601 585
R1146 VSS.n601 VSS.n600 585
R1147 VSS.n2174 VSS.n2173 585
R1148 VSS.n2173 VSS.n2172 585
R1149 VSS.n603 VSS.n602 585
R1150 VSS.n604 VSS.n603 585
R1151 VSS.n2165 VSS.n2164 585
R1152 VSS.n2166 VSS.n2165 585
R1153 VSS.n2163 VSS.n609 585
R1154 VSS.n609 VSS.n608 585
R1155 VSS.n2162 VSS.n2161 585
R1156 VSS.n2161 VSS.n2160 585
R1157 VSS.n611 VSS.n610 585
R1158 VSS.n612 VSS.n611 585
R1159 VSS.n2153 VSS.n2152 585
R1160 VSS.n2154 VSS.n2153 585
R1161 VSS.n2151 VSS.n618 585
R1162 VSS.n618 VSS.n616 585
R1163 VSS.n2150 VSS.n2149 585
R1164 VSS.n2149 VSS.n2148 585
R1165 VSS.n620 VSS.n619 585
R1166 VSS.n621 VSS.n620 585
R1167 VSS.n2141 VSS.n2140 585
R1168 VSS.n2142 VSS.n2141 585
R1169 VSS.n2139 VSS.n626 585
R1170 VSS.n626 VSS.n625 585
R1171 VSS.n2138 VSS.n2137 585
R1172 VSS.n2137 VSS.n2136 585
R1173 VSS.n628 VSS.n627 585
R1174 VSS.n629 VSS.n628 585
R1175 VSS.n2129 VSS.n2128 585
R1176 VSS.n2130 VSS.n2129 585
R1177 VSS.n2127 VSS.n634 585
R1178 VSS.n634 VSS.n633 585
R1179 VSS.n2126 VSS.n2125 585
R1180 VSS.n2125 VSS.n2124 585
R1181 VSS.n636 VSS.n635 585
R1182 VSS.n637 VSS.n636 585
R1183 VSS.n2117 VSS.n2116 585
R1184 VSS.n2118 VSS.n2117 585
R1185 VSS.n2115 VSS.n642 585
R1186 VSS.n2114 VSS.n2113 585
R1187 VSS.n2111 VSS.n643 585
R1188 VSS.n2111 VSS.n641 585
R1189 VSS.n2110 VSS.n2109 585
R1190 VSS.n645 VSS.n640 585
R1191 VSS.n768 VSS.n767 585
R1192 VSS.n2063 VSS.n2062 585
R1193 VSS.n2061 VSS.n779 585
R1194 VSS.n2065 VSS.n779 585
R1195 VSS.n2060 VSS.n2059 585
R1196 VSS.n2058 VSS.n2057 585
R1197 VSS.n2056 VSS.n2055 585
R1198 VSS.n2054 VSS.n2053 585
R1199 VSS.n2052 VSS.n2051 585
R1200 VSS.n2050 VSS.n2049 585
R1201 VSS.n2048 VSS.n2047 585
R1202 VSS.n2046 VSS.n2045 585
R1203 VSS.n2044 VSS.n2043 585
R1204 VSS.n2042 VSS.n2041 585
R1205 VSS.n2040 VSS.n2039 585
R1206 VSS.n2038 VSS.n2037 585
R1207 VSS.n2036 VSS.n2035 585
R1208 VSS.n2034 VSS.n2033 585
R1209 VSS.n2032 VSS.n2031 585
R1210 VSS.n2030 VSS.n2029 585
R1211 VSS.n2028 VSS.n778 585
R1212 VSS.n2065 VSS.n778 585
R1213 VSS.n1461 VSS.n1460 585
R1214 VSS.n1165 VSS.n1129 585
R1215 VSS.n1164 VSS.n1163 585
R1216 VSS.n1162 VSS.n1161 585
R1217 VSS.n1160 VSS.n1159 585
R1218 VSS.n1158 VSS.n1157 585
R1219 VSS.n1156 VSS.n1155 585
R1220 VSS.n1154 VSS.n1153 585
R1221 VSS.n1152 VSS.n1151 585
R1222 VSS.n1150 VSS.n1149 585
R1223 VSS.n1148 VSS.n1147 585
R1224 VSS.n1146 VSS.n1145 585
R1225 VSS.n1144 VSS.n1143 585
R1226 VSS.n1142 VSS.n1141 585
R1227 VSS.n1140 VSS.n1139 585
R1228 VSS.n1138 VSS.n1137 585
R1229 VSS.n1136 VSS.n1135 585
R1230 VSS.n1134 VSS.n1133 585
R1231 VSS.n1132 VSS.n1131 585
R1232 VSS.n1119 VSS.n1118 585
R1233 VSS.n1467 VSS.n1466 585
R1234 VSS.n1466 VSS.n1465 585
R1235 VSS.n1468 VSS.n1117 585
R1236 VSS.n1464 VSS.n1117 585
R1237 VSS.n1470 VSS.n1469 585
R1238 VSS.n1471 VSS.n1470 585
R1239 VSS.n1116 VSS.n1115 585
R1240 VSS.n1472 VSS.n1116 585
R1241 VSS.n1475 VSS.n1474 585
R1242 VSS.n1474 VSS.n1473 585
R1243 VSS.n1476 VSS.n1113 585
R1244 VSS.n1113 VSS.n1111 585
R1245 VSS.n1517 VSS.n1516 585
R1246 VSS.n1518 VSS.n1517 585
R1247 VSS.n1515 VSS.n1114 585
R1248 VSS.n1114 VSS.n1112 585
R1249 VSS.n1514 VSS.n1513 585
R1250 VSS.n1513 VSS.n1512 585
R1251 VSS.n1511 VSS.n1477 585
R1252 VSS.n1511 VSS.n1098 585
R1253 VSS.n1510 VSS.n1509 585
R1254 VSS.n1510 VSS.n1099 585
R1255 VSS.n1508 VSS.n1478 585
R1256 VSS.n1503 VSS.n1478 585
R1257 VSS.n1507 VSS.n1506 585
R1258 VSS.n1506 VSS.n1505 585
R1259 VSS.n1502 VSS.n1479 585
R1260 VSS.n1504 VSS.n1502 585
R1261 VSS.n1501 VSS.n1481 585
R1262 VSS.n1501 VSS.n1500 585
R1263 VSS.n1483 VSS.n1480 585
R1264 VSS.n1499 VSS.n1480 585
R1265 VSS.n1497 VSS.n1496 585
R1266 VSS.n1498 VSS.n1497 585
R1267 VSS.n1495 VSS.n1482 585
R1268 VSS.n1482 VSS.n1016 585
R1269 VSS.n1492 VSS.n1491 585
R1270 VSS.n1491 VSS.n1017 585
R1271 VSS.n1490 VSS.n1485 585
R1272 VSS.n1490 VSS.n1489 585
R1273 VSS.n1487 VSS.n1486 585
R1274 VSS.n1488 VSS.n1487 585
R1275 VSS.n750 VSS.n749 585
R1276 VSS.n752 VSS.n750 585
R1277 VSS.n2100 VSS.n2099 585
R1278 VSS.n2099 VSS.n2098 585
R1279 VSS.n754 VSS.n751 585
R1280 VSS.n2097 VSS.n751 585
R1281 VSS.n2095 VSS.n2094 585
R1282 VSS.n2096 VSS.n2095 585
R1283 VSS.n2093 VSS.n753 585
R1284 VSS.n757 VSS.n753 585
R1285 VSS.n2092 VSS.n2091 585
R1286 VSS.n2091 VSS.n2090 585
R1287 VSS.n756 VSS.n755 585
R1288 VSS.n2089 VSS.n756 585
R1289 VSS.n2087 VSS.n2086 585
R1290 VSS.n2088 VSS.n2087 585
R1291 VSS.n2085 VSS.n758 585
R1292 VSS.n761 VSS.n758 585
R1293 VSS.n2084 VSS.n2083 585
R1294 VSS.n2083 VSS.n2082 585
R1295 VSS.n760 VSS.n759 585
R1296 VSS.n2081 VSS.n760 585
R1297 VSS.n2079 VSS.n2078 585
R1298 VSS.n2080 VSS.n2079 585
R1299 VSS.n2077 VSS.n762 585
R1300 VSS.n765 VSS.n762 585
R1301 VSS.n2076 VSS.n2075 585
R1302 VSS.n2075 VSS.n2074 585
R1303 VSS.n764 VSS.n763 585
R1304 VSS.n2073 VSS.n764 585
R1305 VSS.n2071 VSS.n2070 585
R1306 VSS.n2072 VSS.n2071 585
R1307 VSS.n2069 VSS.n766 585
R1308 VSS.n769 VSS.n766 585
R1309 VSS.n2068 VSS.n2067 585
R1310 VSS.n2067 VSS.n2066 585
R1311 VSS.n1589 VSS.n1588 585
R1312 VSS.n1587 VSS.n1092 585
R1313 VSS.n1586 VSS.n1091 585
R1314 VSS.n1591 VSS.n1091 585
R1315 VSS.n1585 VSS.n1584 585
R1316 VSS.n1583 VSS.n1582 585
R1317 VSS.n1581 VSS.n1580 585
R1318 VSS.n1579 VSS.n1578 585
R1319 VSS.n1577 VSS.n1576 585
R1320 VSS.n1575 VSS.n1574 585
R1321 VSS.n1573 VSS.n1572 585
R1322 VSS.n1571 VSS.n1570 585
R1323 VSS.n1569 VSS.n1568 585
R1324 VSS.n1567 VSS.n1566 585
R1325 VSS.n1565 VSS.n1564 585
R1326 VSS.n1563 VSS.n1562 585
R1327 VSS.n1561 VSS.n1560 585
R1328 VSS.n1559 VSS.n1558 585
R1329 VSS.n1557 VSS.n1556 585
R1330 VSS.n1555 VSS.n1554 585
R1331 VSS.n1553 VSS.n1552 585
R1332 VSS.n1551 VSS.n1550 585
R1333 VSS.n1549 VSS.n1548 585
R1334 VSS.n1547 VSS.n1546 585
R1335 VSS.n1545 VSS.n1095 585
R1336 VSS.n1545 VSS.n1544 585
R1337 VSS.n1525 VSS.n1096 585
R1338 VSS.n1536 VSS.n1096 585
R1339 VSS.n1527 VSS.n1526 585
R1340 VSS.n1528 VSS.n1527 585
R1341 VSS.n1522 VSS.n1107 585
R1342 VSS.n1530 VSS.n1107 585
R1343 VSS.n1521 VSS.n1520 585
R1344 VSS.n1520 VSS.n1519 585
R1345 VSS.n1109 VSS.n1108 585
R1346 VSS.n1309 VSS.n1109 585
R1347 VSS.n1304 VSS.n1303 585
R1348 VSS.n1305 VSS.n1304 585
R1349 VSS.n1302 VSS.n1233 585
R1350 VSS.n1322 VSS.n1233 585
R1351 VSS.n1301 VSS.n1300 585
R1352 VSS.n1300 VSS.n1299 585
R1353 VSS.n1298 VSS.n1225 585
R1354 VSS.n1328 VSS.n1225 585
R1355 VSS.n1297 VSS.n1296 585
R1356 VSS.n1296 VSS.n1224 585
R1357 VSS.n1295 VSS.n1234 585
R1358 VSS.n1295 VSS.n1294 585
R1359 VSS.n1253 VSS.n1235 585
R1360 VSS.n1254 VSS.n1252 585
R1361 VSS.n1256 VSS.n1255 585
R1362 VSS.n1258 VSS.n1249 585
R1363 VSS.n1260 VSS.n1259 585
R1364 VSS.n1261 VSS.n1248 585
R1365 VSS.n1263 VSS.n1262 585
R1366 VSS.n1265 VSS.n1246 585
R1367 VSS.n1267 VSS.n1266 585
R1368 VSS.n1268 VSS.n1245 585
R1369 VSS.n1270 VSS.n1269 585
R1370 VSS.n1272 VSS.n1243 585
R1371 VSS.n1274 VSS.n1273 585
R1372 VSS.n1275 VSS.n1242 585
R1373 VSS.n1277 VSS.n1276 585
R1374 VSS.n1279 VSS.n1240 585
R1375 VSS.n1281 VSS.n1280 585
R1376 VSS.n1282 VSS.n1239 585
R1377 VSS.n1284 VSS.n1283 585
R1378 VSS.n1286 VSS.n1238 585
R1379 VSS.n1287 VSS.n1237 585
R1380 VSS.n1290 VSS.n1289 585
R1381 VSS.n1291 VSS.n1236 585
R1382 VSS.n1236 VSS.n139 585
R1383 VSS.n1293 VSS.n1292 585
R1384 VSS.n1294 VSS.n1293 585
R1385 VSS.n1229 VSS.n1227 585
R1386 VSS.n1227 VSS.n1224 585
R1387 VSS.n1327 VSS.n1326 585
R1388 VSS.n1328 VSS.n1327 585
R1389 VSS.n1325 VSS.n1228 585
R1390 VSS.n1299 VSS.n1228 585
R1391 VSS.n1324 VSS.n1323 585
R1392 VSS.n1323 VSS.n1322 585
R1393 VSS.n1231 VSS.n1230 585
R1394 VSS.n1305 VSS.n1231 585
R1395 VSS.n1308 VSS.n1307 585
R1396 VSS.n1309 VSS.n1308 585
R1397 VSS.n1105 VSS.n1104 585
R1398 VSS.n1519 VSS.n1105 585
R1399 VSS.n1532 VSS.n1531 585
R1400 VSS.n1531 VSS.n1530 585
R1401 VSS.n1533 VSS.n1103 585
R1402 VSS.n1528 VSS.n1103 585
R1403 VSS.n1535 VSS.n1534 585
R1404 VSS.n1536 VSS.n1535 585
R1405 VSS.n1094 VSS.n1093 585
R1406 VSS.n1544 VSS.n1093 585
R1407 VSS.n1865 VSS.n836 585
R1408 VSS.n1864 VSS.n1863 585
R1409 VSS.n1861 VSS.n838 585
R1410 VSS.n1861 VSS.n835 585
R1411 VSS.n1860 VSS.n1859 585
R1412 VSS.n1858 VSS.n1857 585
R1413 VSS.n1856 VSS.n840 585
R1414 VSS.n1854 VSS.n1853 585
R1415 VSS.n1852 VSS.n841 585
R1416 VSS.n1851 VSS.n1850 585
R1417 VSS.n1848 VSS.n842 585
R1418 VSS.n1846 VSS.n1845 585
R1419 VSS.n1842 VSS.n843 585
R1420 VSS.n1841 VSS.n1840 585
R1421 VSS.n1838 VSS.n845 585
R1422 VSS.n1836 VSS.n1835 585
R1423 VSS.n1834 VSS.n846 585
R1424 VSS.n1833 VSS.n1832 585
R1425 VSS.n1830 VSS.n847 585
R1426 VSS.n1828 VSS.n1827 585
R1427 VSS.n1826 VSS.n848 585
R1428 VSS.n1825 VSS.n1824 585
R1429 VSS.n1822 VSS.n849 585
R1430 VSS.n1820 VSS.n1819 585
R1431 VSS.n1818 VSS.n834 585
R1432 VSS.n1868 VSS.n834 585
R1433 VSS.n1817 VSS.n833 585
R1434 VSS.n1869 VSS.n833 585
R1435 VSS.n1816 VSS.n832 585
R1436 VSS.n1870 VSS.n832 585
R1437 VSS.n1815 VSS.n1814 585
R1438 VSS.n1814 VSS.n820 585
R1439 VSS.n1813 VSS.n819 585
R1440 VSS.n2024 VSS.n819 585
R1441 VSS.n1812 VSS.n1811 585
R1442 VSS.n1811 VSS.n782 585
R1443 VSS.n1810 VSS.n826 585
R1444 VSS.n1878 VSS.n826 585
R1445 VSS.n1809 VSS.n1808 585
R1446 VSS.n1808 VSS.n1807 585
R1447 VSS.n1806 VSS.n850 585
R1448 VSS.n1806 VSS.n1805 585
R1449 VSS.n1737 VSS.n851 585
R1450 VSS.n859 VSS.n851 585
R1451 VSS.n1738 VSS.n858 585
R1452 VSS.n1799 VSS.n858 585
R1453 VSS.n1741 VSS.n1739 585
R1454 VSS.n1741 VSS.n1740 585
R1455 VSS.n1743 VSS.n1742 585
R1456 VSS.n1745 VSS.n1744 585
R1457 VSS.n1747 VSS.n1746 585
R1458 VSS.n1749 VSS.n1748 585
R1459 VSS.n1751 VSS.n1750 585
R1460 VSS.n1753 VSS.n1752 585
R1461 VSS.n1755 VSS.n1754 585
R1462 VSS.n1757 VSS.n1756 585
R1463 VSS.n1759 VSS.n1758 585
R1464 VSS.n1761 VSS.n1760 585
R1465 VSS.n1763 VSS.n1762 585
R1466 VSS.n1765 VSS.n1764 585
R1467 VSS.n1767 VSS.n1766 585
R1468 VSS.n1769 VSS.n1768 585
R1469 VSS.n1771 VSS.n1770 585
R1470 VSS.n1773 VSS.n1772 585
R1471 VSS.n1775 VSS.n1774 585
R1472 VSS.n1777 VSS.n1776 585
R1473 VSS.n1779 VSS.n1778 585
R1474 VSS.n1781 VSS.n1780 585
R1475 VSS.n1783 VSS.n1782 585
R1476 VSS.n1784 VSS.n1736 585
R1477 VSS.n1786 VSS.n1785 585
R1478 VSS.n1787 VSS.n1786 585
R1479 VSS.n856 VSS.n855 585
R1480 VSS.n1740 VSS.n856 585
R1481 VSS.n1801 VSS.n1800 585
R1482 VSS.n1800 VSS.n1799 585
R1483 VSS.n1802 VSS.n854 585
R1484 VSS.n859 VSS.n854 585
R1485 VSS.n1804 VSS.n1803 585
R1486 VSS.n1805 VSS.n1804 585
R1487 VSS.n829 VSS.n827 585
R1488 VSS.n1807 VSS.n827 585
R1489 VSS.n1877 VSS.n1876 585
R1490 VSS.n1878 VSS.n1877 585
R1491 VSS.n1875 VSS.n828 585
R1492 VSS.n828 VSS.n782 585
R1493 VSS.n1874 VSS.n821 585
R1494 VSS.n2024 VSS.n821 585
R1495 VSS.n1873 VSS.n1872 585
R1496 VSS.n1872 VSS.n820 585
R1497 VSS.n1871 VSS.n830 585
R1498 VSS.n1871 VSS.n1870 585
R1499 VSS.n837 VSS.n831 585
R1500 VSS.n1869 VSS.n831 585
R1501 VSS.n1867 VSS.n1866 585
R1502 VSS.n1868 VSS.n1867 585
R1503 VSS.n2540 VSS.n2539 585
R1504 VSS.n2538 VSS.n141 585
R1505 VSS.n2537 VSS.n140 585
R1506 VSS.n2542 VSS.n140 585
R1507 VSS.n2536 VSS.n2535 585
R1508 VSS.n2534 VSS.n2533 585
R1509 VSS.n2532 VSS.n2531 585
R1510 VSS.n2530 VSS.n2529 585
R1511 VSS.n2528 VSS.n2527 585
R1512 VSS.n2526 VSS.n2525 585
R1513 VSS.n2524 VSS.n2523 585
R1514 VSS.n2522 VSS.n2521 585
R1515 VSS.n2520 VSS.n2519 585
R1516 VSS.n2518 VSS.n2517 585
R1517 VSS.n2516 VSS.n2515 585
R1518 VSS.n2514 VSS.n2513 585
R1519 VSS.n2512 VSS.n2511 585
R1520 VSS.n2510 VSS.n2509 585
R1521 VSS.n2508 VSS.n2507 585
R1522 VSS.n2506 VSS.n2505 585
R1523 VSS.n2504 VSS.n2503 585
R1524 VSS.n2494 VSS.n2493 585
R1525 VSS.n2496 VSS.n2495 585
R1526 VSS.n2499 VSS.n2498 585
R1527 VSS.n120 VSS.n117 585
R1528 VSS.n2545 VSS.n2544 585
R1529 VSS.n119 VSS.n118 585
R1530 VSS.n2461 VSS.n2460 585
R1531 VSS.n2463 VSS.n2462 585
R1532 VSS.n2465 VSS.n2464 585
R1533 VSS.n2467 VSS.n2466 585
R1534 VSS.n2469 VSS.n2468 585
R1535 VSS.n2471 VSS.n2470 585
R1536 VSS.n2473 VSS.n2472 585
R1537 VSS.n2475 VSS.n2474 585
R1538 VSS.n2477 VSS.n2476 585
R1539 VSS.n2479 VSS.n2478 585
R1540 VSS.n2481 VSS.n2480 585
R1541 VSS.n2483 VSS.n2482 585
R1542 VSS.n2485 VSS.n2484 585
R1543 VSS.n2486 VSS.n147 585
R1544 VSS.n147 VSS.n121 585
R1545 VSS.n2488 VSS.n2487 585
R1546 VSS.n2489 VSS.n2488 585
R1547 VSS.n2459 VSS.n146 585
R1548 VSS.n146 VSS.n145 585
R1549 VSS.n2458 VSS.n2457 585
R1550 VSS.n2457 VSS.n2456 585
R1551 VSS.n149 VSS.n148 585
R1552 VSS.n150 VSS.n149 585
R1553 VSS.n2449 VSS.n2448 585
R1554 VSS.n2450 VSS.n2449 585
R1555 VSS.n2447 VSS.n154 585
R1556 VSS.n158 VSS.n154 585
R1557 VSS.n2446 VSS.n2445 585
R1558 VSS.n2445 VSS.n2444 585
R1559 VSS.n156 VSS.n155 585
R1560 VSS.n157 VSS.n156 585
R1561 VSS.n2437 VSS.n2436 585
R1562 VSS.n2438 VSS.n2437 585
R1563 VSS.n2435 VSS.n162 585
R1564 VSS.n166 VSS.n162 585
R1565 VSS.n2434 VSS.n2433 585
R1566 VSS.n2433 VSS.n2432 585
R1567 VSS.n164 VSS.n163 585
R1568 VSS.n165 VSS.n164 585
R1569 VSS.n2425 VSS.n2424 585
R1570 VSS.n2426 VSS.n2425 585
R1571 VSS.n2423 VSS.n170 585
R1572 VSS.n174 VSS.n170 585
R1573 VSS.n2422 VSS.n2421 585
R1574 VSS.n2421 VSS.n2420 585
R1575 VSS.n172 VSS.n171 585
R1576 VSS.n173 VSS.n172 585
R1577 VSS.n2413 VSS.n2412 585
R1578 VSS.n2414 VSS.n2413 585
R1579 VSS.n2411 VSS.n178 585
R1580 VSS.n182 VSS.n178 585
R1581 VSS.n2410 VSS.n2409 585
R1582 VSS.n2409 VSS.n2408 585
R1583 VSS.n180 VSS.n179 585
R1584 VSS.n181 VSS.n180 585
R1585 VSS.n2401 VSS.n2400 585
R1586 VSS.n2402 VSS.n2401 585
R1587 VSS.n2399 VSS.n186 585
R1588 VSS.n190 VSS.n186 585
R1589 VSS.n2398 VSS.n2397 585
R1590 VSS.n2397 VSS.n2396 585
R1591 VSS.n188 VSS.n187 585
R1592 VSS.n189 VSS.n188 585
R1593 VSS.n2389 VSS.n2388 585
R1594 VSS.n2390 VSS.n2389 585
R1595 VSS.n2387 VSS.n195 585
R1596 VSS.n195 VSS.n194 585
R1597 VSS.n2386 VSS.n2385 585
R1598 VSS.n2385 VSS.n2384 585
R1599 VSS.n197 VSS.n196 585
R1600 VSS.n198 VSS.n197 585
R1601 VSS.n2377 VSS.n2376 585
R1602 VSS.n2378 VSS.n2377 585
R1603 VSS.n2375 VSS.n203 585
R1604 VSS.n203 VSS.n202 585
R1605 VSS.n2374 VSS.n2373 585
R1606 VSS.n2373 VSS.n2372 585
R1607 VSS.n205 VSS.n204 585
R1608 VSS.n206 VSS.n205 585
R1609 VSS.n2365 VSS.n2364 585
R1610 VSS.n2366 VSS.n2365 585
R1611 VSS.n2363 VSS.n211 585
R1612 VSS.n211 VSS.n210 585
R1613 VSS.n2362 VSS.n2361 585
R1614 VSS.n2361 VSS.n2360 585
R1615 VSS.n213 VSS.n212 585
R1616 VSS.n214 VSS.n213 585
R1617 VSS.n2353 VSS.n2352 585
R1618 VSS.n2354 VSS.n2353 585
R1619 VSS.n2351 VSS.n219 585
R1620 VSS.n219 VSS.n218 585
R1621 VSS.n2350 VSS.n2349 585
R1622 VSS.n2349 VSS.n2348 585
R1623 VSS.n221 VSS.n220 585
R1624 VSS.n2341 VSS.n221 585
R1625 VSS.n2340 VSS.n2339 585
R1626 VSS.n2342 VSS.n2340 585
R1627 VSS.n2338 VSS.n226 585
R1628 VSS.n226 VSS.n225 585
R1629 VSS.n2337 VSS.n2336 585
R1630 VSS.n2336 VSS.n2335 585
R1631 VSS.n228 VSS.n227 585
R1632 VSS.n2328 VSS.n228 585
R1633 VSS.n2327 VSS.n2326 585
R1634 VSS.n2329 VSS.n2327 585
R1635 VSS.n2325 VSS.n233 585
R1636 VSS.n233 VSS.n232 585
R1637 VSS.n2324 VSS.n2323 585
R1638 VSS.n2323 VSS.n2322 585
R1639 VSS.n235 VSS.n234 585
R1640 VSS.n2315 VSS.n235 585
R1641 VSS.n2314 VSS.n2313 585
R1642 VSS.n2316 VSS.n2314 585
R1643 VSS.n2312 VSS.n240 585
R1644 VSS.n240 VSS.n239 585
R1645 VSS.n2311 VSS.n2310 585
R1646 VSS.n2310 VSS.n2309 585
R1647 VSS.n242 VSS.n241 585
R1648 VSS.n2302 VSS.n242 585
R1649 VSS.n2301 VSS.n2300 585
R1650 VSS.n2303 VSS.n2301 585
R1651 VSS.n2299 VSS.n247 585
R1652 VSS.n247 VSS.n246 585
R1653 VSS.n2298 VSS.n2297 585
R1654 VSS.n2297 VSS.n2296 585
R1655 VSS.n249 VSS.n248 585
R1656 VSS.n2288 VSS.n249 585
R1657 VSS.n526 VSS.n525 585
R1658 VSS.n2290 VSS.n526 585
R1659 VSS.n524 VSS.n254 585
R1660 VSS.n254 VSS.n253 585
R1661 VSS.n523 VSS.n522 585
R1662 VSS.n522 VSS.n521 585
R1663 VSS.n256 VSS.n255 585
R1664 VSS.n257 VSS.n256 585
R1665 VSS.n514 VSS.n513 585
R1666 VSS.n515 VSS.n514 585
R1667 VSS.n512 VSS.n262 585
R1668 VSS.n511 VSS.n510 585
R1669 VSS.n508 VSS.n263 585
R1670 VSS.n506 VSS.n505 585
R1671 VSS.n504 VSS.n264 585
R1672 VSS.n503 VSS.n502 585
R1673 VSS.n500 VSS.n265 585
R1674 VSS.n498 VSS.n497 585
R1675 VSS.n496 VSS.n266 585
R1676 VSS.n495 VSS.n494 585
R1677 VSS.n492 VSS.n267 585
R1678 VSS.n490 VSS.n489 585
R1679 VSS.n488 VSS.n268 585
R1680 VSS.n487 VSS.n486 585
R1681 VSS.n484 VSS.n269 585
R1682 VSS.n482 VSS.n481 585
R1683 VSS.n271 VSS.n270 585
R1684 VSS.n325 VSS.n324 585
R1685 VSS.n322 VSS.n273 585
R1686 VSS.n320 VSS.n319 585
R1687 VSS.n318 VSS.n274 585
R1688 VSS.n317 VSS.n316 585
R1689 VSS.n314 VSS.n275 585
R1690 VSS.n312 VSS.n311 585
R1691 VSS.n310 VSS.n276 585
R1692 VSS.n309 VSS.n308 585
R1693 VSS.n306 VSS.n277 585
R1694 VSS.n304 VSS.n303 585
R1695 VSS.n302 VSS.n278 585
R1696 VSS.n301 VSS.n300 585
R1697 VSS.n298 VSS.n279 585
R1698 VSS.n296 VSS.n295 585
R1699 VSS.n294 VSS.n280 585
R1700 VSS.n293 VSS.n292 585
R1701 VSS.n290 VSS.n281 585
R1702 VSS.n288 VSS.n287 585
R1703 VSS.n286 VSS.n282 585
R1704 VSS.n285 VSS.n284 585
R1705 VSS.n260 VSS.n259 585
R1706 VSS.n261 VSS.n260 585
R1707 VSS.n517 VSS.n516 585
R1708 VSS.n516 VSS.n515 585
R1709 VSS.n518 VSS.n258 585
R1710 VSS.n258 VSS.n257 585
R1711 VSS.n520 VSS.n519 585
R1712 VSS.n521 VSS.n520 585
R1713 VSS.n252 VSS.n251 585
R1714 VSS.n253 VSS.n252 585
R1715 VSS.n2292 VSS.n2291 585
R1716 VSS.n2291 VSS.n2290 585
R1717 VSS.n2293 VSS.n250 585
R1718 VSS.n2288 VSS.n250 585
R1719 VSS.n2295 VSS.n2294 585
R1720 VSS.n2296 VSS.n2295 585
R1721 VSS.n245 VSS.n244 585
R1722 VSS.n246 VSS.n245 585
R1723 VSS.n2305 VSS.n2304 585
R1724 VSS.n2304 VSS.n2303 585
R1725 VSS.n2306 VSS.n243 585
R1726 VSS.n2302 VSS.n243 585
R1727 VSS.n2308 VSS.n2307 585
R1728 VSS.n2309 VSS.n2308 585
R1729 VSS.n238 VSS.n237 585
R1730 VSS.n239 VSS.n238 585
R1731 VSS.n2318 VSS.n2317 585
R1732 VSS.n2317 VSS.n2316 585
R1733 VSS.n2319 VSS.n236 585
R1734 VSS.n2315 VSS.n236 585
R1735 VSS.n2321 VSS.n2320 585
R1736 VSS.n2322 VSS.n2321 585
R1737 VSS.n231 VSS.n230 585
R1738 VSS.n232 VSS.n231 585
R1739 VSS.n2331 VSS.n2330 585
R1740 VSS.n2330 VSS.n2329 585
R1741 VSS.n2332 VSS.n229 585
R1742 VSS.n2328 VSS.n229 585
R1743 VSS.n2334 VSS.n2333 585
R1744 VSS.n2335 VSS.n2334 585
R1745 VSS.n224 VSS.n223 585
R1746 VSS.n225 VSS.n224 585
R1747 VSS.n2344 VSS.n2343 585
R1748 VSS.n2343 VSS.n2342 585
R1749 VSS.n2345 VSS.n222 585
R1750 VSS.n2341 VSS.n222 585
R1751 VSS.n2347 VSS.n2346 585
R1752 VSS.n2348 VSS.n2347 585
R1753 VSS.n217 VSS.n216 585
R1754 VSS.n218 VSS.n217 585
R1755 VSS.n2356 VSS.n2355 585
R1756 VSS.n2355 VSS.n2354 585
R1757 VSS.n2357 VSS.n215 585
R1758 VSS.n215 VSS.n214 585
R1759 VSS.n2359 VSS.n2358 585
R1760 VSS.n2360 VSS.n2359 585
R1761 VSS.n209 VSS.n208 585
R1762 VSS.n210 VSS.n209 585
R1763 VSS.n2368 VSS.n2367 585
R1764 VSS.n2367 VSS.n2366 585
R1765 VSS.n2369 VSS.n207 585
R1766 VSS.n207 VSS.n206 585
R1767 VSS.n2371 VSS.n2370 585
R1768 VSS.n2372 VSS.n2371 585
R1769 VSS.n201 VSS.n200 585
R1770 VSS.n202 VSS.n201 585
R1771 VSS.n2380 VSS.n2379 585
R1772 VSS.n2379 VSS.n2378 585
R1773 VSS.n2381 VSS.n199 585
R1774 VSS.n199 VSS.n198 585
R1775 VSS.n2383 VSS.n2382 585
R1776 VSS.n2384 VSS.n2383 585
R1777 VSS.n193 VSS.n192 585
R1778 VSS.n194 VSS.n193 585
R1779 VSS.n2392 VSS.n2391 585
R1780 VSS.n2391 VSS.n2390 585
R1781 VSS.n2393 VSS.n191 585
R1782 VSS.n191 VSS.n189 585
R1783 VSS.n2395 VSS.n2394 585
R1784 VSS.n2396 VSS.n2395 585
R1785 VSS.n185 VSS.n184 585
R1786 VSS.n190 VSS.n185 585
R1787 VSS.n2404 VSS.n2403 585
R1788 VSS.n2403 VSS.n2402 585
R1789 VSS.n2405 VSS.n183 585
R1790 VSS.n183 VSS.n181 585
R1791 VSS.n2407 VSS.n2406 585
R1792 VSS.n2408 VSS.n2407 585
R1793 VSS.n177 VSS.n176 585
R1794 VSS.n182 VSS.n177 585
R1795 VSS.n2416 VSS.n2415 585
R1796 VSS.n2415 VSS.n2414 585
R1797 VSS.n2417 VSS.n175 585
R1798 VSS.n175 VSS.n173 585
R1799 VSS.n2419 VSS.n2418 585
R1800 VSS.n2420 VSS.n2419 585
R1801 VSS.n169 VSS.n168 585
R1802 VSS.n174 VSS.n169 585
R1803 VSS.n2428 VSS.n2427 585
R1804 VSS.n2427 VSS.n2426 585
R1805 VSS.n2429 VSS.n167 585
R1806 VSS.n167 VSS.n165 585
R1807 VSS.n2431 VSS.n2430 585
R1808 VSS.n2432 VSS.n2431 585
R1809 VSS.n161 VSS.n160 585
R1810 VSS.n166 VSS.n161 585
R1811 VSS.n2440 VSS.n2439 585
R1812 VSS.n2439 VSS.n2438 585
R1813 VSS.n2441 VSS.n159 585
R1814 VSS.n159 VSS.n157 585
R1815 VSS.n2443 VSS.n2442 585
R1816 VSS.n2444 VSS.n2443 585
R1817 VSS.n153 VSS.n152 585
R1818 VSS.n158 VSS.n153 585
R1819 VSS.n2452 VSS.n2451 585
R1820 VSS.n2451 VSS.n2450 585
R1821 VSS.n2453 VSS.n151 585
R1822 VSS.n151 VSS.n150 585
R1823 VSS.n2455 VSS.n2454 585
R1824 VSS.n2456 VSS.n2455 585
R1825 VSS.n144 VSS.n143 585
R1826 VSS.n145 VSS.n144 585
R1827 VSS.n2491 VSS.n2490 585
R1828 VSS.n2490 VSS.n2489 585
R1829 VSS.n2492 VSS.n142 585
R1830 VSS.n142 VSS.n121 585
R1831 VSS.n2027 VSS.n2026 585
R1832 VSS.n781 VSS.n780 585
R1833 VSS.n2023 VSS.n2022 585
R1834 VSS.n2024 VSS.n2023 585
R1835 VSS.n2021 VSS.n822 585
R1836 VSS.n2020 VSS.n2019 585
R1837 VSS.n2018 VSS.n2017 585
R1838 VSS.n2016 VSS.n2015 585
R1839 VSS.n2014 VSS.n2013 585
R1840 VSS.n2012 VSS.n2011 585
R1841 VSS.n2010 VSS.n2009 585
R1842 VSS.n2008 VSS.n2007 585
R1843 VSS.n2006 VSS.n2005 585
R1844 VSS.n2004 VSS.n2003 585
R1845 VSS.n2002 VSS.n2001 585
R1846 VSS.n2000 VSS.n1999 585
R1847 VSS.n1998 VSS.n1997 585
R1848 VSS.n1996 VSS.n1995 585
R1849 VSS.n1994 VSS.n1993 585
R1850 VSS.n1992 VSS.n1991 585
R1851 VSS.n1990 VSS.n1989 585
R1852 VSS.n1988 VSS.n1987 585
R1853 VSS.n1986 VSS.n1985 585
R1854 VSS.n1984 VSS.n1983 585
R1855 VSS.n1982 VSS.n1981 585
R1856 VSS.n1980 VSS.n1979 585
R1857 VSS.n1978 VSS.n1977 585
R1858 VSS.n1976 VSS.n1975 585
R1859 VSS.n1974 VSS.n1973 585
R1860 VSS.n1972 VSS.n1971 585
R1861 VSS.n1970 VSS.n1969 585
R1862 VSS.n1968 VSS.n1967 585
R1863 VSS.n1966 VSS.n1965 585
R1864 VSS.n1964 VSS.n1963 585
R1865 VSS.n1962 VSS.n1961 585
R1866 VSS.n1960 VSS.n1959 585
R1867 VSS.n1958 VSS.n1957 585
R1868 VSS.n1956 VSS.n1955 585
R1869 VSS.n1954 VSS.n1953 585
R1870 VSS.n1952 VSS.n1951 585
R1871 VSS.n1950 VSS.n1949 585
R1872 VSS.n1948 VSS.n1947 585
R1873 VSS.n1946 VSS.n1945 585
R1874 VSS.n1944 VSS.n1943 585
R1875 VSS.n1942 VSS.n1941 585
R1876 VSS.n1940 VSS.n1939 585
R1877 VSS.n1938 VSS.n1937 585
R1878 VSS.n1936 VSS.n1935 585
R1879 VSS.n1934 VSS.n1933 585
R1880 VSS.n1932 VSS.n1931 585
R1881 VSS.n1930 VSS.n1929 585
R1882 VSS.n1928 VSS.n1927 585
R1883 VSS.n1926 VSS.n1925 585
R1884 VSS.n1924 VSS.n1923 585
R1885 VSS.n1922 VSS.n1921 585
R1886 VSS.n1920 VSS.n1919 585
R1887 VSS.n1918 VSS.n1917 585
R1888 VSS.n1916 VSS.n1915 585
R1889 VSS.n1914 VSS.n1913 585
R1890 VSS.n1912 VSS.n1911 585
R1891 VSS.n1910 VSS.n1909 585
R1892 VSS.n1908 VSS.n1907 585
R1893 VSS.n1906 VSS.n1905 585
R1894 VSS.n1904 VSS.n1903 585
R1895 VSS.n1902 VSS.n1901 585
R1896 VSS.n1900 VSS.n1899 585
R1897 VSS.n1898 VSS.n1897 585
R1898 VSS.n1896 VSS.n1895 585
R1899 VSS.n1894 VSS.n1893 585
R1900 VSS.n1892 VSS.n1891 585
R1901 VSS.n1890 VSS.n1889 585
R1902 VSS.n1888 VSS.n1887 585
R1903 VSS.n1886 VSS.n1885 585
R1904 VSS.n1884 VSS.n1883 585
R1905 VSS.n1882 VSS.n818 585
R1906 VSS.n2024 VSS.n818 585
R1907 VSS.n1881 VSS.n1880 585
R1908 VSS.n1880 VSS.n1879 585
R1909 VSS.n824 VSS.n823 585
R1910 VSS.n825 VSS.n824 585
R1911 VSS.n1794 VSS.n1793 585
R1912 VSS.n1793 VSS.n853 585
R1913 VSS.n1795 VSS.n861 585
R1914 VSS.n861 VSS.n852 585
R1915 VSS.n1797 VSS.n1796 585
R1916 VSS.n1798 VSS.n1797 585
R1917 VSS.n1792 VSS.n860 585
R1918 VSS.n860 VSS.n857 585
R1919 VSS.n1791 VSS.n1790 585
R1920 VSS.n1790 VSS.n1789 585
R1921 VSS.n863 VSS.n862 585
R1922 VSS.n1788 VSS.n863 585
R1923 VSS.n1723 VSS.n1722 585
R1924 VSS.n1724 VSS.n1723 585
R1925 VSS.n1721 VSS.n865 585
R1926 VSS.n865 VSS.n864 585
R1927 VSS.n1720 VSS.n1719 585
R1928 VSS.n1719 VSS.n1718 585
R1929 VSS.n867 VSS.n866 585
R1930 VSS.n868 VSS.n867 585
R1931 VSS.n1668 VSS.n1667 585
R1932 VSS.n1669 VSS.n1668 585
R1933 VSS.n1666 VSS.n887 585
R1934 VSS.n887 VSS.n886 585
R1935 VSS.n1665 VSS.n1664 585
R1936 VSS.n1664 VSS.n1663 585
R1937 VSS.n889 VSS.n888 585
R1938 VSS.n1654 VSS.n889 585
R1939 VSS.n1628 VSS.n1627 585
R1940 VSS.n1628 VSS.n896 585
R1941 VSS.n1632 VSS.n1631 585
R1942 VSS.n1631 VSS.n1630 585
R1943 VSS.n1633 VSS.n909 585
R1944 VSS.n909 VSS.n901 585
R1945 VSS.n1635 VSS.n1634 585
R1946 VSS.n1636 VSS.n1635 585
R1947 VSS.n910 VSS.n908 585
R1948 VSS.n908 VSS.n905 585
R1949 VSS.n1619 VSS.n1618 585
R1950 VSS.n1618 VSS.n1617 585
R1951 VSS.n1014 VSS.n1013 585
R1952 VSS.n1022 VSS.n1014 585
R1953 VSS.n1597 VSS.n1077 585
R1954 VSS.n1077 VSS.n1021 585
R1955 VSS.n1599 VSS.n1598 585
R1956 VSS.n1600 VSS.n1599 585
R1957 VSS.n1596 VSS.n1076 585
R1958 VSS.n1592 VSS.n1076 585
R1959 VSS.n1595 VSS.n1594 585
R1960 VSS.n1594 VSS.n1593 585
R1961 VSS.n1079 VSS.n1078 585
R1962 VSS.n1080 VSS.n1079 585
R1963 VSS.n1542 VSS.n1541 585
R1964 VSS.n1543 VSS.n1542 585
R1965 VSS.n1540 VSS.n1100 585
R1966 VSS.n1100 VSS.n1097 585
R1967 VSS.n1539 VSS.n1538 585
R1968 VSS.n1538 VSS.n1537 585
R1969 VSS.n1102 VSS.n1101 585
R1970 VSS.n1529 VSS.n1102 585
R1971 VSS.n1315 VSS.n1314 585
R1972 VSS.n1315 VSS.n1106 585
R1973 VSS.n1317 VSS.n1316 585
R1974 VSS.n1316 VSS.n1110 585
R1975 VSS.n1318 VSS.n1311 585
R1976 VSS.n1311 VSS.n1310 585
R1977 VSS.n1320 VSS.n1319 585
R1978 VSS.n1321 VSS.n1320 585
R1979 VSS.n1313 VSS.n1306 585
R1980 VSS.n1306 VSS.n1232 585
R1981 VSS.n1312 VSS.n1223 585
R1982 VSS.n1226 VSS.n1223 585
R1983 VSS.n1330 VSS.n1221 585
R1984 VSS.n1330 VSS.n1329 585
R1985 VSS.n1332 VSS.n1331 585
R1986 VSS.n1333 VSS.n1220 585
R1987 VSS.n1335 VSS.n1334 585
R1988 VSS.n1337 VSS.n1218 585
R1989 VSS.n1339 VSS.n1338 585
R1990 VSS.n1340 VSS.n1217 585
R1991 VSS.n1342 VSS.n1341 585
R1992 VSS.n1344 VSS.n1215 585
R1993 VSS.n1346 VSS.n1345 585
R1994 VSS.n1347 VSS.n1214 585
R1995 VSS.n1349 VSS.n1348 585
R1996 VSS.n1351 VSS.n1212 585
R1997 VSS.n1353 VSS.n1352 585
R1998 VSS.n1354 VSS.n1211 585
R1999 VSS.n1356 VSS.n1355 585
R2000 VSS.n1358 VSS.n1209 585
R2001 VSS.n1360 VSS.n1359 585
R2002 VSS.n1361 VSS.n1208 585
R2003 VSS.n1363 VSS.n1362 585
R2004 VSS.n1365 VSS.n1206 585
R2005 VSS.n1367 VSS.n1366 585
R2006 VSS.n1368 VSS.n1205 585
R2007 VSS.n1370 VSS.n1369 585
R2008 VSS.n1372 VSS.n1203 585
R2009 VSS.n1374 VSS.n1373 585
R2010 VSS.n1375 VSS.n1202 585
R2011 VSS.n1377 VSS.n1376 585
R2012 VSS.n1379 VSS.n1200 585
R2013 VSS.n1381 VSS.n1380 585
R2014 VSS.n1382 VSS.n1199 585
R2015 VSS.n1384 VSS.n1383 585
R2016 VSS.n1386 VSS.n1197 585
R2017 VSS.n1388 VSS.n1387 585
R2018 VSS.n1389 VSS.n1196 585
R2019 VSS.n1391 VSS.n1390 585
R2020 VSS.n1393 VSS.n1194 585
R2021 VSS.n1395 VSS.n1394 585
R2022 VSS.n1396 VSS.n1193 585
R2023 VSS.n1398 VSS.n1397 585
R2024 VSS.n1400 VSS.n1191 585
R2025 VSS.n1402 VSS.n1401 585
R2026 VSS.n1403 VSS.n1190 585
R2027 VSS.n1405 VSS.n1404 585
R2028 VSS.n1407 VSS.n1188 585
R2029 VSS.n1409 VSS.n1408 585
R2030 VSS.n1410 VSS.n1187 585
R2031 VSS.n1412 VSS.n1411 585
R2032 VSS.n1414 VSS.n1185 585
R2033 VSS.n1416 VSS.n1415 585
R2034 VSS.n1417 VSS.n1184 585
R2035 VSS.n1419 VSS.n1418 585
R2036 VSS.n1421 VSS.n1182 585
R2037 VSS.n1423 VSS.n1422 585
R2038 VSS.n1424 VSS.n1181 585
R2039 VSS.n1426 VSS.n1425 585
R2040 VSS.n1428 VSS.n1179 585
R2041 VSS.n1430 VSS.n1429 585
R2042 VSS.n1431 VSS.n1178 585
R2043 VSS.n1433 VSS.n1432 585
R2044 VSS.n1435 VSS.n1176 585
R2045 VSS.n1437 VSS.n1436 585
R2046 VSS.n1438 VSS.n1175 585
R2047 VSS.n1440 VSS.n1439 585
R2048 VSS.n1442 VSS.n1173 585
R2049 VSS.n1444 VSS.n1443 585
R2050 VSS.n1445 VSS.n1172 585
R2051 VSS.n1447 VSS.n1446 585
R2052 VSS.n1449 VSS.n1170 585
R2053 VSS.n1451 VSS.n1450 585
R2054 VSS.n1452 VSS.n1169 585
R2055 VSS.n1454 VSS.n1453 585
R2056 VSS.n1456 VSS.n1166 585
R2057 VSS.n1458 VSS.n1457 585
R2058 VSS.n1459 VSS.n1130 585
R2059 VSS.n1020 VSS.n1019 585
R2060 VSS.n1601 VSS.n1020 585
R2061 VSS.n1074 VSS.n1073 585
R2062 VSS.n1072 VSS.n1037 585
R2063 VSS.n1071 VSS.n1070 585
R2064 VSS.n1069 VSS.n1068 585
R2065 VSS.n1067 VSS.n1066 585
R2066 VSS.n1065 VSS.n1064 585
R2067 VSS.n1063 VSS.n1062 585
R2068 VSS.n1061 VSS.n1060 585
R2069 VSS.n1059 VSS.n1058 585
R2070 VSS.n1057 VSS.n1056 585
R2071 VSS.n1055 VSS.n1054 585
R2072 VSS.n1053 VSS.n1052 585
R2073 VSS.n1051 VSS.n1050 585
R2074 VSS.n1049 VSS.n1048 585
R2075 VSS.n1047 VSS.n1046 585
R2076 VSS.n1045 VSS.n1044 585
R2077 VSS.n1043 VSS.n1042 585
R2078 VSS.n1041 VSS.n1040 585
R2079 VSS.n1039 VSS.n1038 585
R2080 VSS.n1027 VSS.n1026 585
R2081 VSS.n1604 VSS.n1603 585
R2082 VSS.n1605 VSS.n1023 585
R2083 VSS.n1608 VSS.n1607 585
R2084 VSS.n1609 VSS.n1608 585
R2085 VSS.n1606 VSS.n1025 585
R2086 VSS.n1025 VSS.n1024 585
R2087 VSS.n904 VSS.n903 585
R2088 VSS.n1616 VSS.n904 585
R2089 VSS.n1639 VSS.n1638 585
R2090 VSS.n1638 VSS.n1637 585
R2091 VSS.n1640 VSS.n902 585
R2092 VSS.n907 VSS.n902 585
R2093 VSS.n1642 VSS.n1641 585
R2094 VSS.n1643 VSS.n1642 585
R2095 VSS.n895 VSS.n894 585
R2096 VSS.n1629 VSS.n895 585
R2097 VSS.n1657 VSS.n1656 585
R2098 VSS.n1656 VSS.n1655 585
R2099 VSS.n1658 VSS.n892 585
R2100 VSS.n892 VSS.n890 585
R2101 VSS.n1661 VSS.n1660 585
R2102 VSS.n1662 VSS.n1661 585
R2103 VSS.n1659 VSS.n893 585
R2104 VSS.n893 VSS.n885 585
R2105 VSS.n882 VSS.n881 585
R2106 VSS.n1670 VSS.n881 585
R2107 VSS.n1715 VSS.n1714 585
R2108 VSS.n1713 VSS.n880 585
R2109 VSS.n1712 VSS.n879 585
R2110 VSS.n1717 VSS.n879 585
R2111 VSS.n1711 VSS.n1710 585
R2112 VSS.n1709 VSS.n1708 585
R2113 VSS.n1707 VSS.n1706 585
R2114 VSS.n1705 VSS.n1704 585
R2115 VSS.n1703 VSS.n1702 585
R2116 VSS.n1701 VSS.n1700 585
R2117 VSS.n1699 VSS.n1698 585
R2118 VSS.n1697 VSS.n1696 585
R2119 VSS.n1695 VSS.n1694 585
R2120 VSS.n1693 VSS.n1692 585
R2121 VSS.n1691 VSS.n1690 585
R2122 VSS.n1689 VSS.n1688 585
R2123 VSS.n1687 VSS.n1686 585
R2124 VSS.n1685 VSS.n1684 585
R2125 VSS.n1683 VSS.n1682 585
R2126 VSS.n1681 VSS.n1680 585
R2127 VSS.n1679 VSS.n1678 585
R2128 VSS.n1677 VSS.n1676 585
R2129 VSS.n1675 VSS.n1674 585
R2130 VSS.n1673 VSS.n1672 585
R2131 VSS.n1671 VSS.n883 585
R2132 VSS.n1671 VSS.n1670 585
R2133 VSS.n1647 VSS.n884 585
R2134 VSS.n885 VSS.n884 585
R2135 VSS.n1648 VSS.n891 585
R2136 VSS.n1662 VSS.n891 585
R2137 VSS.n1650 VSS.n898 585
R2138 VSS.n898 VSS.n890 585
R2139 VSS.n1653 VSS.n1652 585
R2140 VSS.n1655 VSS.n1653 585
R2141 VSS.n1646 VSS.n897 585
R2142 VSS.n1629 VSS.n897 585
R2143 VSS.n1645 VSS.n1644 585
R2144 VSS.n1644 VSS.n1643 585
R2145 VSS.n900 VSS.n899 585
R2146 VSS.n907 VSS.n900 585
R2147 VSS.n1613 VSS.n906 585
R2148 VSS.n1637 VSS.n906 585
R2149 VSS.n1615 VSS.n1614 585
R2150 VSS.n1616 VSS.n1615 585
R2151 VSS.n1612 VSS.n1018 585
R2152 VSS.n1024 VSS.n1018 585
R2153 VSS.n1611 VSS.n1610 585
R2154 VSS.n1610 VSS.n1609 585
R2155 VSS.n516 VSS.n258 394
R2156 VSS.n520 VSS.n258 394
R2157 VSS.n520 VSS.n252 394
R2158 VSS.n2291 VSS.n252 394
R2159 VSS.n2291 VSS.n250 394
R2160 VSS.n2295 VSS.n250 394
R2161 VSS.n2295 VSS.n245 394
R2162 VSS.n2304 VSS.n245 394
R2163 VSS.n2304 VSS.n243 394
R2164 VSS.n2308 VSS.n243 394
R2165 VSS.n2308 VSS.n238 394
R2166 VSS.n2317 VSS.n238 394
R2167 VSS.n2317 VSS.n236 394
R2168 VSS.n2321 VSS.n236 394
R2169 VSS.n2321 VSS.n231 394
R2170 VSS.n2330 VSS.n231 394
R2171 VSS.n2330 VSS.n229 394
R2172 VSS.n2334 VSS.n229 394
R2173 VSS.n2334 VSS.n224 394
R2174 VSS.n2343 VSS.n224 394
R2175 VSS.n2343 VSS.n222 394
R2176 VSS.n2347 VSS.n222 394
R2177 VSS.n2347 VSS.n217 394
R2178 VSS.n2355 VSS.n217 394
R2179 VSS.n2355 VSS.n215 394
R2180 VSS.n2359 VSS.n215 394
R2181 VSS.n2359 VSS.n209 394
R2182 VSS.n2367 VSS.n209 394
R2183 VSS.n2367 VSS.n207 394
R2184 VSS.n2371 VSS.n207 394
R2185 VSS.n2371 VSS.n201 394
R2186 VSS.n2379 VSS.n201 394
R2187 VSS.n2379 VSS.n199 394
R2188 VSS.n2383 VSS.n199 394
R2189 VSS.n2383 VSS.n193 394
R2190 VSS.n2391 VSS.n193 394
R2191 VSS.n2391 VSS.n191 394
R2192 VSS.n2395 VSS.n191 394
R2193 VSS.n2395 VSS.n185 394
R2194 VSS.n2403 VSS.n185 394
R2195 VSS.n2403 VSS.n183 394
R2196 VSS.n2407 VSS.n183 394
R2197 VSS.n2407 VSS.n177 394
R2198 VSS.n2415 VSS.n177 394
R2199 VSS.n2415 VSS.n175 394
R2200 VSS.n2419 VSS.n175 394
R2201 VSS.n2419 VSS.n169 394
R2202 VSS.n2427 VSS.n169 394
R2203 VSS.n2427 VSS.n167 394
R2204 VSS.n2431 VSS.n167 394
R2205 VSS.n2431 VSS.n161 394
R2206 VSS.n2439 VSS.n161 394
R2207 VSS.n2439 VSS.n159 394
R2208 VSS.n2443 VSS.n159 394
R2209 VSS.n2443 VSS.n153 394
R2210 VSS.n2451 VSS.n153 394
R2211 VSS.n2451 VSS.n151 394
R2212 VSS.n2455 VSS.n151 394
R2213 VSS.n2455 VSS.n144 394
R2214 VSS.n2490 VSS.n144 394
R2215 VSS.n2490 VSS.n142 394
R2216 VSS.n284 VSS.n260 394
R2217 VSS.n288 VSS.n282 394
R2218 VSS.n292 VSS.n290 394
R2219 VSS.n296 VSS.n280 394
R2220 VSS.n300 VSS.n298 394
R2221 VSS.n304 VSS.n278 394
R2222 VSS.n308 VSS.n306 394
R2223 VSS.n312 VSS.n276 394
R2224 VSS.n316 VSS.n314 394
R2225 VSS.n320 VSS.n274 394
R2226 VSS.n324 VSS.n322 394
R2227 VSS.n482 VSS.n270 394
R2228 VSS.n486 VSS.n484 394
R2229 VSS.n490 VSS.n268 394
R2230 VSS.n494 VSS.n492 394
R2231 VSS.n498 VSS.n266 394
R2232 VSS.n502 VSS.n500 394
R2233 VSS.n506 VSS.n264 394
R2234 VSS.n510 VSS.n508 394
R2235 VSS.n514 VSS.n256 394
R2236 VSS.n522 VSS.n256 394
R2237 VSS.n522 VSS.n254 394
R2238 VSS.n526 VSS.n254 394
R2239 VSS.n526 VSS.n249 394
R2240 VSS.n2297 VSS.n249 394
R2241 VSS.n2297 VSS.n247 394
R2242 VSS.n2301 VSS.n247 394
R2243 VSS.n2301 VSS.n242 394
R2244 VSS.n2310 VSS.n242 394
R2245 VSS.n2310 VSS.n240 394
R2246 VSS.n2314 VSS.n240 394
R2247 VSS.n2314 VSS.n235 394
R2248 VSS.n2323 VSS.n235 394
R2249 VSS.n2323 VSS.n233 394
R2250 VSS.n2327 VSS.n233 394
R2251 VSS.n2327 VSS.n228 394
R2252 VSS.n2336 VSS.n228 394
R2253 VSS.n2336 VSS.n226 394
R2254 VSS.n2340 VSS.n226 394
R2255 VSS.n2340 VSS.n221 394
R2256 VSS.n2349 VSS.n221 394
R2257 VSS.n2349 VSS.n219 394
R2258 VSS.n2353 VSS.n219 394
R2259 VSS.n2353 VSS.n213 394
R2260 VSS.n2361 VSS.n213 394
R2261 VSS.n2361 VSS.n211 394
R2262 VSS.n2365 VSS.n211 394
R2263 VSS.n2365 VSS.n205 394
R2264 VSS.n2373 VSS.n205 394
R2265 VSS.n2373 VSS.n203 394
R2266 VSS.n2377 VSS.n203 394
R2267 VSS.n2377 VSS.n197 394
R2268 VSS.n2385 VSS.n197 394
R2269 VSS.n2385 VSS.n195 394
R2270 VSS.n2389 VSS.n195 394
R2271 VSS.n2389 VSS.n188 394
R2272 VSS.n2397 VSS.n188 394
R2273 VSS.n2397 VSS.n186 394
R2274 VSS.n2401 VSS.n186 394
R2275 VSS.n2401 VSS.n180 394
R2276 VSS.n2409 VSS.n180 394
R2277 VSS.n2409 VSS.n178 394
R2278 VSS.n2413 VSS.n178 394
R2279 VSS.n2413 VSS.n172 394
R2280 VSS.n2421 VSS.n172 394
R2281 VSS.n2421 VSS.n170 394
R2282 VSS.n2425 VSS.n170 394
R2283 VSS.n2425 VSS.n164 394
R2284 VSS.n2433 VSS.n164 394
R2285 VSS.n2433 VSS.n162 394
R2286 VSS.n2437 VSS.n162 394
R2287 VSS.n2437 VSS.n156 394
R2288 VSS.n2445 VSS.n156 394
R2289 VSS.n2445 VSS.n154 394
R2290 VSS.n2449 VSS.n154 394
R2291 VSS.n2449 VSS.n149 394
R2292 VSS.n2457 VSS.n149 394
R2293 VSS.n2457 VSS.n146 394
R2294 VSS.n2488 VSS.n146 394
R2295 VSS.n2488 VSS.n147 394
R2296 VSS.n141 VSS.n140 394
R2297 VSS.n2535 VSS.n140 394
R2298 VSS.n2533 VSS.n2532 394
R2299 VSS.n2529 VSS.n2528 394
R2300 VSS.n2525 VSS.n2524 394
R2301 VSS.n2521 VSS.n2520 394
R2302 VSS.n2517 VSS.n2516 394
R2303 VSS.n2513 VSS.n2512 394
R2304 VSS.n2509 VSS.n2508 394
R2305 VSS.n2505 VSS.n2504 394
R2306 VSS.n2495 VSS.n2494 394
R2307 VSS.n2498 VSS.n120 394
R2308 VSS.n2544 VSS.n119 394
R2309 VSS.n2462 VSS.n2461 394
R2310 VSS.n2466 VSS.n2465 394
R2311 VSS.n2470 VSS.n2469 394
R2312 VSS.n2474 VSS.n2473 394
R2313 VSS.n2478 VSS.n2477 394
R2314 VSS.n2482 VSS.n2481 394
R2315 VSS.n1800 VSS.n856 394
R2316 VSS.n1800 VSS.n854 394
R2317 VSS.n1804 VSS.n854 394
R2318 VSS.n1804 VSS.n827 394
R2319 VSS.n1877 VSS.n827 394
R2320 VSS.n1877 VSS.n828 394
R2321 VSS.n828 VSS.n821 394
R2322 VSS.n1872 VSS.n821 394
R2323 VSS.n1872 VSS.n1871 394
R2324 VSS.n1871 VSS.n831 394
R2325 VSS.n1867 VSS.n831 394
R2326 VSS.n1786 VSS.n1736 394
R2327 VSS.n1782 VSS.n1781 394
R2328 VSS.n1778 VSS.n1777 394
R2329 VSS.n1774 VSS.n1773 394
R2330 VSS.n1770 VSS.n1769 394
R2331 VSS.n1766 VSS.n1765 394
R2332 VSS.n1762 VSS.n1761 394
R2333 VSS.n1758 VSS.n1757 394
R2334 VSS.n1754 VSS.n1753 394
R2335 VSS.n1750 VSS.n1749 394
R2336 VSS.n1746 VSS.n1745 394
R2337 VSS.n1741 VSS.n858 394
R2338 VSS.n858 VSS.n851 394
R2339 VSS.n1806 VSS.n851 394
R2340 VSS.n1808 VSS.n1806 394
R2341 VSS.n1808 VSS.n826 394
R2342 VSS.n1811 VSS.n826 394
R2343 VSS.n1811 VSS.n819 394
R2344 VSS.n1814 VSS.n819 394
R2345 VSS.n1814 VSS.n832 394
R2346 VSS.n833 VSS.n832 394
R2347 VSS.n834 VSS.n833 394
R2348 VSS.n1863 VSS.n1861 394
R2349 VSS.n1861 VSS.n1860 394
R2350 VSS.n1857 VSS.n1856 394
R2351 VSS.n1854 VSS.n841 394
R2352 VSS.n1850 VSS.n1848 394
R2353 VSS.n1846 VSS.n843 394
R2354 VSS.n1840 VSS.n1838 394
R2355 VSS.n1836 VSS.n846 394
R2356 VSS.n1832 VSS.n1830 394
R2357 VSS.n1828 VSS.n848 394
R2358 VSS.n1824 VSS.n1822 394
R2359 VSS.n1293 VSS.n1227 394
R2360 VSS.n1327 VSS.n1227 394
R2361 VSS.n1327 VSS.n1228 394
R2362 VSS.n1323 VSS.n1228 394
R2363 VSS.n1323 VSS.n1231 394
R2364 VSS.n1308 VSS.n1231 394
R2365 VSS.n1308 VSS.n1105 394
R2366 VSS.n1531 VSS.n1105 394
R2367 VSS.n1531 VSS.n1103 394
R2368 VSS.n1535 VSS.n1103 394
R2369 VSS.n1535 VSS.n1093 394
R2370 VSS.n1289 VSS.n1236 394
R2371 VSS.n1287 VSS.n1286 394
R2372 VSS.n1284 VSS.n1239 394
R2373 VSS.n1280 VSS.n1279 394
R2374 VSS.n1277 VSS.n1242 394
R2375 VSS.n1273 VSS.n1272 394
R2376 VSS.n1270 VSS.n1245 394
R2377 VSS.n1266 VSS.n1265 394
R2378 VSS.n1263 VSS.n1248 394
R2379 VSS.n1259 VSS.n1258 394
R2380 VSS.n1256 VSS.n1252 394
R2381 VSS.n1296 VSS.n1295 394
R2382 VSS.n1296 VSS.n1225 394
R2383 VSS.n1300 VSS.n1225 394
R2384 VSS.n1300 VSS.n1233 394
R2385 VSS.n1304 VSS.n1233 394
R2386 VSS.n1304 VSS.n1109 394
R2387 VSS.n1520 VSS.n1109 394
R2388 VSS.n1520 VSS.n1107 394
R2389 VSS.n1527 VSS.n1107 394
R2390 VSS.n1527 VSS.n1096 394
R2391 VSS.n1545 VSS.n1096 394
R2392 VSS.n1092 VSS.n1091 394
R2393 VSS.n1584 VSS.n1091 394
R2394 VSS.n1582 VSS.n1581 394
R2395 VSS.n1578 VSS.n1577 394
R2396 VSS.n1574 VSS.n1573 394
R2397 VSS.n1570 VSS.n1569 394
R2398 VSS.n1566 VSS.n1565 394
R2399 VSS.n1562 VSS.n1561 394
R2400 VSS.n1558 VSS.n1557 394
R2401 VSS.n1554 VSS.n1553 394
R2402 VSS.n1550 VSS.n1549 394
R2403 VSS.n1466 VSS.n1117 394
R2404 VSS.n1470 VSS.n1117 394
R2405 VSS.n1470 VSS.n1116 394
R2406 VSS.n1474 VSS.n1116 394
R2407 VSS.n1474 VSS.n1113 394
R2408 VSS.n1517 VSS.n1113 394
R2409 VSS.n1517 VSS.n1114 394
R2410 VSS.n1513 VSS.n1114 394
R2411 VSS.n1513 VSS.n1511 394
R2412 VSS.n1511 VSS.n1510 394
R2413 VSS.n1510 VSS.n1478 394
R2414 VSS.n1506 VSS.n1478 394
R2415 VSS.n1506 VSS.n1502 394
R2416 VSS.n1502 VSS.n1501 394
R2417 VSS.n1501 VSS.n1480 394
R2418 VSS.n1497 VSS.n1480 394
R2419 VSS.n1497 VSS.n1482 394
R2420 VSS.n1491 VSS.n1482 394
R2421 VSS.n1491 VSS.n1490 394
R2422 VSS.n1490 VSS.n1487 394
R2423 VSS.n1487 VSS.n750 394
R2424 VSS.n2099 VSS.n750 394
R2425 VSS.n2099 VSS.n751 394
R2426 VSS.n2095 VSS.n751 394
R2427 VSS.n2095 VSS.n753 394
R2428 VSS.n2091 VSS.n753 394
R2429 VSS.n2091 VSS.n756 394
R2430 VSS.n2087 VSS.n756 394
R2431 VSS.n2087 VSS.n758 394
R2432 VSS.n2083 VSS.n758 394
R2433 VSS.n2083 VSS.n760 394
R2434 VSS.n2079 VSS.n760 394
R2435 VSS.n2079 VSS.n762 394
R2436 VSS.n2075 VSS.n762 394
R2437 VSS.n2075 VSS.n764 394
R2438 VSS.n2071 VSS.n764 394
R2439 VSS.n2071 VSS.n766 394
R2440 VSS.n2067 VSS.n766 394
R2441 VSS.n1133 VSS.n1132 394
R2442 VSS.n1137 VSS.n1136 394
R2443 VSS.n1141 VSS.n1140 394
R2444 VSS.n1145 VSS.n1144 394
R2445 VSS.n1149 VSS.n1148 394
R2446 VSS.n1153 VSS.n1152 394
R2447 VSS.n1157 VSS.n1156 394
R2448 VSS.n1161 VSS.n1160 394
R2449 VSS.n1163 VSS.n1129 394
R2450 VSS.n1461 VSS.n1130 394
R2451 VSS.n1457 VSS.n1456 394
R2452 VSS.n1454 VSS.n1169 394
R2453 VSS.n1450 VSS.n1449 394
R2454 VSS.n1447 VSS.n1172 394
R2455 VSS.n1443 VSS.n1442 394
R2456 VSS.n1440 VSS.n1175 394
R2457 VSS.n1436 VSS.n1435 394
R2458 VSS.n1433 VSS.n1178 394
R2459 VSS.n1429 VSS.n1428 394
R2460 VSS.n1426 VSS.n1181 394
R2461 VSS.n1422 VSS.n1421 394
R2462 VSS.n1419 VSS.n1184 394
R2463 VSS.n1415 VSS.n1414 394
R2464 VSS.n1412 VSS.n1187 394
R2465 VSS.n1408 VSS.n1407 394
R2466 VSS.n1405 VSS.n1190 394
R2467 VSS.n1401 VSS.n1400 394
R2468 VSS.n1398 VSS.n1193 394
R2469 VSS.n1394 VSS.n1393 394
R2470 VSS.n1391 VSS.n1196 394
R2471 VSS.n1387 VSS.n1386 394
R2472 VSS.n1384 VSS.n1199 394
R2473 VSS.n1380 VSS.n1379 394
R2474 VSS.n1377 VSS.n1202 394
R2475 VSS.n1373 VSS.n1372 394
R2476 VSS.n1370 VSS.n1205 394
R2477 VSS.n1366 VSS.n1365 394
R2478 VSS.n1363 VSS.n1208 394
R2479 VSS.n1359 VSS.n1358 394
R2480 VSS.n1356 VSS.n1211 394
R2481 VSS.n1352 VSS.n1351 394
R2482 VSS.n1349 VSS.n1214 394
R2483 VSS.n1345 VSS.n1344 394
R2484 VSS.n1342 VSS.n1217 394
R2485 VSS.n1338 VSS.n1337 394
R2486 VSS.n1335 VSS.n1220 394
R2487 VSS.n1330 VSS.n1223 394
R2488 VSS.n1306 VSS.n1223 394
R2489 VSS.n1320 VSS.n1306 394
R2490 VSS.n1320 VSS.n1311 394
R2491 VSS.n1316 VSS.n1311 394
R2492 VSS.n1316 VSS.n1315 394
R2493 VSS.n1315 VSS.n1102 394
R2494 VSS.n1538 VSS.n1102 394
R2495 VSS.n1538 VSS.n1100 394
R2496 VSS.n1542 VSS.n1100 394
R2497 VSS.n1542 VSS.n1079 394
R2498 VSS.n1594 VSS.n1079 394
R2499 VSS.n1594 VSS.n1076 394
R2500 VSS.n1599 VSS.n1076 394
R2501 VSS.n1599 VSS.n1077 394
R2502 VSS.n1077 VSS.n1014 394
R2503 VSS.n1618 VSS.n1014 394
R2504 VSS.n1618 VSS.n908 394
R2505 VSS.n1635 VSS.n908 394
R2506 VSS.n1635 VSS.n909 394
R2507 VSS.n1631 VSS.n909 394
R2508 VSS.n1631 VSS.n1628 394
R2509 VSS.n1628 VSS.n889 394
R2510 VSS.n1664 VSS.n889 394
R2511 VSS.n1664 VSS.n887 394
R2512 VSS.n1668 VSS.n887 394
R2513 VSS.n1668 VSS.n867 394
R2514 VSS.n1719 VSS.n867 394
R2515 VSS.n1719 VSS.n865 394
R2516 VSS.n1723 VSS.n865 394
R2517 VSS.n1723 VSS.n863 394
R2518 VSS.n1790 VSS.n863 394
R2519 VSS.n1790 VSS.n860 394
R2520 VSS.n1797 VSS.n860 394
R2521 VSS.n1797 VSS.n861 394
R2522 VSS.n1793 VSS.n861 394
R2523 VSS.n1793 VSS.n824 394
R2524 VSS.n1880 VSS.n824 394
R2525 VSS.n2063 VSS.n779 394
R2526 VSS.n2059 VSS.n779 394
R2527 VSS.n2057 VSS.n2056 394
R2528 VSS.n2053 VSS.n2052 394
R2529 VSS.n2049 VSS.n2048 394
R2530 VSS.n2045 VSS.n2044 394
R2531 VSS.n2041 VSS.n2040 394
R2532 VSS.n2037 VSS.n2036 394
R2533 VSS.n2033 VSS.n2032 394
R2534 VSS.n2029 VSS.n778 394
R2535 VSS.n2026 VSS.n778 394
R2536 VSS.n2023 VSS.n781 394
R2537 VSS.n2019 VSS.n2018 394
R2538 VSS.n2015 VSS.n2014 394
R2539 VSS.n2011 VSS.n2010 394
R2540 VSS.n2007 VSS.n2006 394
R2541 VSS.n2003 VSS.n2002 394
R2542 VSS.n1999 VSS.n1998 394
R2543 VSS.n1995 VSS.n1994 394
R2544 VSS.n1991 VSS.n1990 394
R2545 VSS.n1987 VSS.n1986 394
R2546 VSS.n1983 VSS.n1982 394
R2547 VSS.n1979 VSS.n1978 394
R2548 VSS.n1971 VSS.n1970 394
R2549 VSS.n1967 VSS.n1966 394
R2550 VSS.n1963 VSS.n1962 394
R2551 VSS.n1959 VSS.n1958 394
R2552 VSS.n1955 VSS.n1954 394
R2553 VSS.n1951 VSS.n1950 394
R2554 VSS.n1947 VSS.n1946 394
R2555 VSS.n1943 VSS.n1942 394
R2556 VSS.n1939 VSS.n1938 394
R2557 VSS.n1935 VSS.n1934 394
R2558 VSS.n1931 VSS.n1930 394
R2559 VSS.n1923 VSS.n1922 394
R2560 VSS.n1919 VSS.n1918 394
R2561 VSS.n1915 VSS.n1914 394
R2562 VSS.n1911 VSS.n1910 394
R2563 VSS.n1907 VSS.n1906 394
R2564 VSS.n1903 VSS.n1902 394
R2565 VSS.n1899 VSS.n1898 394
R2566 VSS.n1895 VSS.n1894 394
R2567 VSS.n1891 VSS.n1890 394
R2568 VSS.n1887 VSS.n1886 394
R2569 VSS.n1883 VSS.n818 394
R2570 VSS.n2113 VSS.n2111 394
R2571 VSS.n2111 VSS.n2110 394
R2572 VSS.n2117 VSS.n636 394
R2573 VSS.n2125 VSS.n636 394
R2574 VSS.n2125 VSS.n634 394
R2575 VSS.n2129 VSS.n634 394
R2576 VSS.n2129 VSS.n628 394
R2577 VSS.n2137 VSS.n628 394
R2578 VSS.n2137 VSS.n626 394
R2579 VSS.n2141 VSS.n626 394
R2580 VSS.n2141 VSS.n620 394
R2581 VSS.n2149 VSS.n620 394
R2582 VSS.n2149 VSS.n618 394
R2583 VSS.n2153 VSS.n618 394
R2584 VSS.n2153 VSS.n611 394
R2585 VSS.n2161 VSS.n611 394
R2586 VSS.n2161 VSS.n609 394
R2587 VSS.n2165 VSS.n609 394
R2588 VSS.n2165 VSS.n603 394
R2589 VSS.n2173 VSS.n603 394
R2590 VSS.n2173 VSS.n601 394
R2591 VSS.n2177 VSS.n601 394
R2592 VSS.n2177 VSS.n595 394
R2593 VSS.n2185 VSS.n595 394
R2594 VSS.n2185 VSS.n593 394
R2595 VSS.n2189 VSS.n593 394
R2596 VSS.n2189 VSS.n587 394
R2597 VSS.n2197 VSS.n587 394
R2598 VSS.n2197 VSS.n585 394
R2599 VSS.n2201 VSS.n585 394
R2600 VSS.n2201 VSS.n579 394
R2601 VSS.n2209 VSS.n579 394
R2602 VSS.n2209 VSS.n577 394
R2603 VSS.n2213 VSS.n577 394
R2604 VSS.n2213 VSS.n571 394
R2605 VSS.n2221 VSS.n571 394
R2606 VSS.n2221 VSS.n569 394
R2607 VSS.n2225 VSS.n569 394
R2608 VSS.n2225 VSS.n563 394
R2609 VSS.n2233 VSS.n563 394
R2610 VSS.n2233 VSS.n561 394
R2611 VSS.n2237 VSS.n561 394
R2612 VSS.n2237 VSS.n555 394
R2613 VSS.n2245 VSS.n555 394
R2614 VSS.n2245 VSS.n553 394
R2615 VSS.n2249 VSS.n553 394
R2616 VSS.n2249 VSS.n547 394
R2617 VSS.n2257 VSS.n547 394
R2618 VSS.n2257 VSS.n545 394
R2619 VSS.n2261 VSS.n545 394
R2620 VSS.n2261 VSS.n539 394
R2621 VSS.n2270 VSS.n539 394
R2622 VSS.n2270 VSS.n537 394
R2623 VSS.n2274 VSS.n537 394
R2624 VSS.n2274 VSS.n530 394
R2625 VSS.n2286 VSS.n531 394
R2626 VSS.n2282 VSS.n2281 394
R2627 VSS.n2119 VSS.n638 394
R2628 VSS.n2123 VSS.n638 394
R2629 VSS.n2123 VSS.n632 394
R2630 VSS.n2131 VSS.n632 394
R2631 VSS.n2131 VSS.n630 394
R2632 VSS.n2135 VSS.n630 394
R2633 VSS.n2135 VSS.n624 394
R2634 VSS.n2143 VSS.n624 394
R2635 VSS.n2143 VSS.n622 394
R2636 VSS.n2147 VSS.n622 394
R2637 VSS.n2147 VSS.n615 394
R2638 VSS.n2155 VSS.n615 394
R2639 VSS.n2155 VSS.n613 394
R2640 VSS.n2159 VSS.n613 394
R2641 VSS.n2159 VSS.n607 394
R2642 VSS.n2167 VSS.n607 394
R2643 VSS.n2167 VSS.n605 394
R2644 VSS.n2171 VSS.n605 394
R2645 VSS.n2171 VSS.n599 394
R2646 VSS.n2179 VSS.n599 394
R2647 VSS.n2179 VSS.n597 394
R2648 VSS.n2183 VSS.n597 394
R2649 VSS.n2183 VSS.n591 394
R2650 VSS.n2191 VSS.n591 394
R2651 VSS.n2191 VSS.n589 394
R2652 VSS.n2195 VSS.n589 394
R2653 VSS.n2195 VSS.n583 394
R2654 VSS.n2203 VSS.n583 394
R2655 VSS.n2203 VSS.n581 394
R2656 VSS.n2207 VSS.n581 394
R2657 VSS.n2207 VSS.n575 394
R2658 VSS.n2215 VSS.n575 394
R2659 VSS.n2215 VSS.n573 394
R2660 VSS.n2219 VSS.n573 394
R2661 VSS.n2219 VSS.n567 394
R2662 VSS.n2227 VSS.n567 394
R2663 VSS.n2227 VSS.n565 394
R2664 VSS.n2231 VSS.n565 394
R2665 VSS.n2231 VSS.n559 394
R2666 VSS.n2239 VSS.n559 394
R2667 VSS.n2239 VSS.n557 394
R2668 VSS.n2243 VSS.n557 394
R2669 VSS.n2243 VSS.n551 394
R2670 VSS.n2251 VSS.n551 394
R2671 VSS.n2251 VSS.n549 394
R2672 VSS.n2255 VSS.n549 394
R2673 VSS.n2255 VSS.n543 394
R2674 VSS.n2263 VSS.n543 394
R2675 VSS.n2263 VSS.n541 394
R2676 VSS.n2268 VSS.n541 394
R2677 VSS.n2268 VSS.n534 394
R2678 VSS.n2276 VSS.n534 394
R2679 VSS.n2277 VSS.n2276 394
R2680 VSS.n1608 VSS.n1025 394
R2681 VSS.n1025 VSS.n904 394
R2682 VSS.n1638 VSS.n904 394
R2683 VSS.n1638 VSS.n902 394
R2684 VSS.n1642 VSS.n902 394
R2685 VSS.n1642 VSS.n895 394
R2686 VSS.n1656 VSS.n895 394
R2687 VSS.n1656 VSS.n892 394
R2688 VSS.n1661 VSS.n892 394
R2689 VSS.n1661 VSS.n893 394
R2690 VSS.n893 VSS.n881 394
R2691 VSS.n880 VSS.n879 394
R2692 VSS.n1710 VSS.n879 394
R2693 VSS.n1708 VSS.n1707 394
R2694 VSS.n1704 VSS.n1703 394
R2695 VSS.n1700 VSS.n1699 394
R2696 VSS.n1696 VSS.n1695 394
R2697 VSS.n1692 VSS.n1691 394
R2698 VSS.n1688 VSS.n1687 394
R2699 VSS.n1684 VSS.n1683 394
R2700 VSS.n1680 VSS.n1679 394
R2701 VSS.n1676 VSS.n1675 394
R2702 VSS.n1610 VSS.n1018 394
R2703 VSS.n1615 VSS.n1018 394
R2704 VSS.n1615 VSS.n906 394
R2705 VSS.n906 VSS.n900 394
R2706 VSS.n1644 VSS.n900 394
R2707 VSS.n1644 VSS.n897 394
R2708 VSS.n1653 VSS.n897 394
R2709 VSS.n1653 VSS.n898 394
R2710 VSS.n898 VSS.n891 394
R2711 VSS.n891 VSS.n884 394
R2712 VSS.n1671 VSS.n884 394
R2713 VSS.n1603 VSS.n1027 394
R2714 VSS.n1040 VSS.n1039 394
R2715 VSS.n1044 VSS.n1043 394
R2716 VSS.n1048 VSS.n1047 394
R2717 VSS.n1052 VSS.n1051 394
R2718 VSS.n1056 VSS.n1055 394
R2719 VSS.n1060 VSS.n1059 394
R2720 VSS.n1064 VSS.n1063 394
R2721 VSS.n1068 VSS.n1067 394
R2722 VSS.n1070 VSS.n1037 394
R2723 VSS.n1074 VSS.n1020 394
R2724 VSS.n2289 VSS.n2287 326.82
R2725 VSS.n112 VSS.n111 325.69
R2726 VSS.n57 VSS.n52 325.69
R2727 VSS.n1455 VSS.n1454 269.089
R2728 VSS.n1456 VSS.n1455 269.089
R2729 VSS.n2542 VSS.n139 261
R2730 VSS.n1001 VSS.t22 259.341
R2731 VSS.n918 VSS.t28 259.341
R2732 VSS.n738 VSS.t121 259.341
R2733 VSS.n655 VSS.t18 259.341
R2734 VSS.n1000 VSS.t145 258.99
R2735 VSS.n999 VSS.t102 258.99
R2736 VSS.n998 VSS.t47 258.99
R2737 VSS.n911 VSS.t108 258.99
R2738 VSS.n912 VSS.t110 258.99
R2739 VSS.n915 VSS.t171 258.99
R2740 VSS.n916 VSS.t10 258.99
R2741 VSS.n917 VSS.t20 258.99
R2742 VSS.n737 VSS.t115 258.99
R2743 VSS.n736 VSS.t100 258.99
R2744 VSS.n735 VSS.t44 258.99
R2745 VSS.n648 VSS.t165 258.99
R2746 VSS.n649 VSS.t129 258.99
R2747 VSS.n652 VSS.t147 258.99
R2748 VSS.n653 VSS.t106 258.99
R2749 VSS.n654 VSS.t51 258.99
R2750 VSS.n996 VSS.n995 253.042
R2751 VSS.n932 VSS.n929 253.042
R2752 VSS.n730 VSS.n700 253.042
R2753 VSS.n670 VSS.n669 253.042
R2754 VSS.n2287 VSS.n528 218.815
R2755 VSS.n2287 VSS.n529 218.815
R2756 VSS.n2112 VSS.n641 218.815
R2757 VSS.n644 VSS.n641 218.815
R2758 VSS.n2065 VSS.n2064 218.815
R2759 VSS.n2065 VSS.n770 218.815
R2760 VSS.n2065 VSS.n771 218.815
R2761 VSS.n2065 VSS.n772 218.815
R2762 VSS.n2065 VSS.n773 218.815
R2763 VSS.n2065 VSS.n774 218.815
R2764 VSS.n2065 VSS.n775 218.815
R2765 VSS.n2065 VSS.n776 218.815
R2766 VSS.n2065 VSS.n777 218.815
R2767 VSS.n1463 VSS.n1462 218.815
R2768 VSS.n1463 VSS.n1128 218.815
R2769 VSS.n1463 VSS.n1127 218.815
R2770 VSS.n1463 VSS.n1126 218.815
R2771 VSS.n1463 VSS.n1125 218.815
R2772 VSS.n1463 VSS.n1124 218.815
R2773 VSS.n1463 VSS.n1123 218.815
R2774 VSS.n1463 VSS.n1122 218.815
R2775 VSS.n1463 VSS.n1121 218.815
R2776 VSS.n1463 VSS.n1120 218.815
R2777 VSS.n1591 VSS.n1590 218.815
R2778 VSS.n1591 VSS.n1081 218.815
R2779 VSS.n1591 VSS.n1082 218.815
R2780 VSS.n1591 VSS.n1083 218.815
R2781 VSS.n1591 VSS.n1084 218.815
R2782 VSS.n1591 VSS.n1085 218.815
R2783 VSS.n1591 VSS.n1086 218.815
R2784 VSS.n1591 VSS.n1087 218.815
R2785 VSS.n1591 VSS.n1088 218.815
R2786 VSS.n1591 VSS.n1089 218.815
R2787 VSS.n1591 VSS.n1090 218.815
R2788 VSS.n1251 VSS.n139 218.815
R2789 VSS.n1257 VSS.n139 218.815
R2790 VSS.n1250 VSS.n139 218.815
R2791 VSS.n1264 VSS.n139 218.815
R2792 VSS.n1247 VSS.n139 218.815
R2793 VSS.n1271 VSS.n139 218.815
R2794 VSS.n1244 VSS.n139 218.815
R2795 VSS.n1278 VSS.n139 218.815
R2796 VSS.n1241 VSS.n139 218.815
R2797 VSS.n1285 VSS.n139 218.815
R2798 VSS.n1288 VSS.n139 218.815
R2799 VSS.n1862 VSS.n835 218.815
R2800 VSS.n839 VSS.n835 218.815
R2801 VSS.n1855 VSS.n835 218.815
R2802 VSS.n1849 VSS.n835 218.815
R2803 VSS.n1847 VSS.n835 218.815
R2804 VSS.n1839 VSS.n835 218.815
R2805 VSS.n1837 VSS.n835 218.815
R2806 VSS.n1831 VSS.n835 218.815
R2807 VSS.n1829 VSS.n835 218.815
R2808 VSS.n1823 VSS.n835 218.815
R2809 VSS.n1821 VSS.n835 218.815
R2810 VSS.n1787 VSS.n1725 218.815
R2811 VSS.n1787 VSS.n1726 218.815
R2812 VSS.n1787 VSS.n1727 218.815
R2813 VSS.n1787 VSS.n1728 218.815
R2814 VSS.n1787 VSS.n1729 218.815
R2815 VSS.n1787 VSS.n1730 218.815
R2816 VSS.n1787 VSS.n1731 218.815
R2817 VSS.n1787 VSS.n1732 218.815
R2818 VSS.n1787 VSS.n1733 218.815
R2819 VSS.n1787 VSS.n1734 218.815
R2820 VSS.n1787 VSS.n1735 218.815
R2821 VSS.n2542 VSS.n2541 218.815
R2822 VSS.n2542 VSS.n122 218.815
R2823 VSS.n2542 VSS.n123 218.815
R2824 VSS.n2542 VSS.n124 218.815
R2825 VSS.n2542 VSS.n125 218.815
R2826 VSS.n2542 VSS.n126 218.815
R2827 VSS.n2542 VSS.n127 218.815
R2828 VSS.n2542 VSS.n128 218.815
R2829 VSS.n2542 VSS.n129 218.815
R2830 VSS.n2542 VSS.n130 218.815
R2831 VSS.n2542 VSS.n131 218.815
R2832 VSS.n2543 VSS.n2542 218.815
R2833 VSS.n2542 VSS.n132 218.815
R2834 VSS.n2542 VSS.n133 218.815
R2835 VSS.n2542 VSS.n134 218.815
R2836 VSS.n2542 VSS.n135 218.815
R2837 VSS.n2542 VSS.n136 218.815
R2838 VSS.n2542 VSS.n137 218.815
R2839 VSS.n2542 VSS.n138 218.815
R2840 VSS.n509 VSS.n261 218.815
R2841 VSS.n507 VSS.n261 218.815
R2842 VSS.n501 VSS.n261 218.815
R2843 VSS.n499 VSS.n261 218.815
R2844 VSS.n493 VSS.n261 218.815
R2845 VSS.n491 VSS.n261 218.815
R2846 VSS.n485 VSS.n261 218.815
R2847 VSS.n483 VSS.n261 218.815
R2848 VSS.n323 VSS.n261 218.815
R2849 VSS.n321 VSS.n261 218.815
R2850 VSS.n315 VSS.n261 218.815
R2851 VSS.n313 VSS.n261 218.815
R2852 VSS.n307 VSS.n261 218.815
R2853 VSS.n305 VSS.n261 218.815
R2854 VSS.n299 VSS.n261 218.815
R2855 VSS.n297 VSS.n261 218.815
R2856 VSS.n291 VSS.n261 218.815
R2857 VSS.n289 VSS.n261 218.815
R2858 VSS.n283 VSS.n261 218.815
R2859 VSS.n2025 VSS.n2024 218.815
R2860 VSS.n2024 VSS.n783 218.815
R2861 VSS.n2024 VSS.n784 218.815
R2862 VSS.n2024 VSS.n785 218.815
R2863 VSS.n2024 VSS.n786 218.815
R2864 VSS.n2024 VSS.n787 218.815
R2865 VSS.n2024 VSS.n788 218.815
R2866 VSS.n2024 VSS.n789 218.815
R2867 VSS.n2024 VSS.n790 218.815
R2868 VSS.n2024 VSS.n791 218.815
R2869 VSS.n2024 VSS.n792 218.815
R2870 VSS.n2024 VSS.n793 218.815
R2871 VSS.n2024 VSS.n794 218.815
R2872 VSS.n2024 VSS.n795 218.815
R2873 VSS.n2024 VSS.n796 218.815
R2874 VSS.n2024 VSS.n797 218.815
R2875 VSS.n2024 VSS.n798 218.815
R2876 VSS.n2024 VSS.n799 218.815
R2877 VSS.n2024 VSS.n800 218.815
R2878 VSS.n2024 VSS.n801 218.815
R2879 VSS.n2024 VSS.n802 218.815
R2880 VSS.n2024 VSS.n803 218.815
R2881 VSS.n2024 VSS.n804 218.815
R2882 VSS.n2024 VSS.n805 218.815
R2883 VSS.n2024 VSS.n806 218.815
R2884 VSS.n2024 VSS.n807 218.815
R2885 VSS.n2024 VSS.n808 218.815
R2886 VSS.n2024 VSS.n809 218.815
R2887 VSS.n2024 VSS.n810 218.815
R2888 VSS.n2024 VSS.n811 218.815
R2889 VSS.n2024 VSS.n812 218.815
R2890 VSS.n2024 VSS.n813 218.815
R2891 VSS.n2024 VSS.n814 218.815
R2892 VSS.n2024 VSS.n815 218.815
R2893 VSS.n2024 VSS.n816 218.815
R2894 VSS.n2024 VSS.n817 218.815
R2895 VSS.n1222 VSS.n1168 218.815
R2896 VSS.n1336 VSS.n1168 218.815
R2897 VSS.n1219 VSS.n1168 218.815
R2898 VSS.n1343 VSS.n1168 218.815
R2899 VSS.n1216 VSS.n1168 218.815
R2900 VSS.n1350 VSS.n1168 218.815
R2901 VSS.n1213 VSS.n1168 218.815
R2902 VSS.n1357 VSS.n1168 218.815
R2903 VSS.n1210 VSS.n1168 218.815
R2904 VSS.n1364 VSS.n1168 218.815
R2905 VSS.n1207 VSS.n1168 218.815
R2906 VSS.n1204 VSS.n1168 218.815
R2907 VSS.n1378 VSS.n1168 218.815
R2908 VSS.n1201 VSS.n1168 218.815
R2909 VSS.n1385 VSS.n1168 218.815
R2910 VSS.n1198 VSS.n1168 218.815
R2911 VSS.n1392 VSS.n1168 218.815
R2912 VSS.n1195 VSS.n1168 218.815
R2913 VSS.n1399 VSS.n1168 218.815
R2914 VSS.n1192 VSS.n1168 218.815
R2915 VSS.n1406 VSS.n1168 218.815
R2916 VSS.n1189 VSS.n1168 218.815
R2917 VSS.n1186 VSS.n1168 218.815
R2918 VSS.n1420 VSS.n1168 218.815
R2919 VSS.n1183 VSS.n1168 218.815
R2920 VSS.n1427 VSS.n1168 218.815
R2921 VSS.n1180 VSS.n1168 218.815
R2922 VSS.n1434 VSS.n1168 218.815
R2923 VSS.n1177 VSS.n1168 218.815
R2924 VSS.n1441 VSS.n1168 218.815
R2925 VSS.n1174 VSS.n1168 218.815
R2926 VSS.n1448 VSS.n1168 218.815
R2927 VSS.n1171 VSS.n1168 218.815
R2928 VSS.n1168 VSS.n1167 218.815
R2929 VSS.n1601 VSS.n1075 218.815
R2930 VSS.n1601 VSS.n1036 218.815
R2931 VSS.n1601 VSS.n1035 218.815
R2932 VSS.n1601 VSS.n1034 218.815
R2933 VSS.n1601 VSS.n1033 218.815
R2934 VSS.n1601 VSS.n1032 218.815
R2935 VSS.n1601 VSS.n1031 218.815
R2936 VSS.n1601 VSS.n1030 218.815
R2937 VSS.n1601 VSS.n1029 218.815
R2938 VSS.n1601 VSS.n1028 218.815
R2939 VSS.n1602 VSS.n1601 218.815
R2940 VSS.n1717 VSS.n1716 218.815
R2941 VSS.n1717 VSS.n869 218.815
R2942 VSS.n1717 VSS.n870 218.815
R2943 VSS.n1717 VSS.n871 218.815
R2944 VSS.n1717 VSS.n872 218.815
R2945 VSS.n1717 VSS.n873 218.815
R2946 VSS.n1717 VSS.n874 218.815
R2947 VSS.n1717 VSS.n875 218.815
R2948 VSS.n1717 VSS.n876 218.815
R2949 VSS.n1717 VSS.n877 218.815
R2950 VSS.n1717 VSS.n878 218.815
R2951 VSS.n2118 VSS.n641 204.464
R2952 VSS.n2287 VSS.n527 204.464
R2953 VSS.n1413 VSS.n1412 198.87
R2954 VSS.n1371 VSS.n1370 198.87
R2955 VSS.n1372 VSS.n1371 198.87
R2956 VSS.n1414 VSS.n1413 198.87
R2957 VSS.n1371 VSS.n1168 193.066
R2958 VSS.n1413 VSS.n1168 193.066
R2959 VSS.n369 VSS.n368 185
R2960 VSS.n369 VSS.n341 185
R2961 VSS.n371 VSS.n370 185
R2962 VSS.n370 VSS.n339 185
R2963 VSS.n353 VSS.n345 185
R2964 VSS.n353 VSS.n344 185
R2965 VSS.n354 VSS.n353 185
R2966 VSS.n474 VSS.n473 185
R2967 VSS.n473 VSS.n457 185
R2968 VSS.n472 VSS.n471 185
R2969 VSS.n472 VSS.n459 185
R2970 VSS.n451 VSS.n443 185
R2971 VSS.n451 VSS.n442 185
R2972 VSS.n452 VSS.n451 185
R2973 VSS.n428 VSS.n427 185
R2974 VSS.n428 VSS.n335 185
R2975 VSS.n428 VSS.n334 185
R2976 VSS.n428 VSS.n332 185
R2977 VSS.n428 VSS.n331 185
R2978 VSS.n428 VSS.n330 185
R2979 VSS.n29 VSS.n11 185
R2980 VSS.n29 VSS.n10 185
R2981 VSS.n29 VSS.n9 185
R2982 VSS.n29 VSS.n8 185
R2983 VSS.n29 VSS.n7 185
R2984 VSS.n29 VSS.n6 185
R2985 VSS.n29 VSS.n5 185
R2986 VSS.n111 VSS.n110 185
R2987 VSS.n88 VSS.n87 185
R2988 VSS.n105 VSS.n104 185
R2989 VSS.n99 VSS.n98 185
R2990 VSS.n99 VSS.n91 185
R2991 VSS.n71 VSS.n70 185
R2992 VSS.n70 VSS.n69 185
R2993 VSS.n57 VSS.n56 185
R2994 VSS.n59 VSS.n58 185
R2995 VSS.n61 VSS.n49 185
R2996 VSS.n974 VSS.n973 185
R2997 VSS.n979 VSS.n978 185
R2998 VSS.n981 VSS.n980 185
R2999 VSS.n970 VSS.n969 185
R3000 VSS.n987 VSS.n986 185
R3001 VSS.n989 VSS.n988 185
R3002 VSS.n966 VSS.n965 185
R3003 VSS.n995 VSS.n994 185
R3004 VSS.n954 VSS.n953 185
R3005 VSS.n922 VSS.n921 185
R3006 VSS.n948 VSS.n947 185
R3007 VSS.n946 VSS.n945 185
R3008 VSS.n926 VSS.n925 185
R3009 VSS.n940 VSS.n939 185
R3010 VSS.n938 VSS.n937 185
R3011 VSS.n930 VSS.n929 185
R3012 VSS.n731 VSS.n730 185
R3013 VSS.n729 VSS.n728 185
R3014 VSS.n704 VSS.n703 185
R3015 VSS.n723 VSS.n722 185
R3016 VSS.n721 VSS.n720 185
R3017 VSS.n708 VSS.n707 185
R3018 VSS.n715 VSS.n714 185
R3019 VSS.n713 VSS.n712 185
R3020 VSS.n671 VSS.n670 185
R3021 VSS.n665 VSS.n664 185
R3022 VSS.n677 VSS.n676 185
R3023 VSS.n679 VSS.n678 185
R3024 VSS.n661 VSS.n660 185
R3025 VSS.n686 VSS.n685 185
R3026 VSS.n688 VSS.n687 185
R3027 VSS.n690 VSS.n657 185
R3028 VSS.n975 VSS.t24 178.418
R3029 VSS.t29 VSS.n920 178.418
R3030 VSS.n711 VSS.t123 178.418
R3031 VSS.t19 VSS.n691 178.418
R3032 VSS.t128 VSS.n103 175.332
R3033 VSS.t156 VSS.n62 175.332
R3034 VSS.n387 VSS.t68 165.607
R3035 VSS.n32 VSS.t15 165.607
R3036 VSS.n399 VSS.t135 165.032
R3037 VSS.n42 VSS.t131 165.032
R3038 VSS.n41 VSS.t167 165.032
R3039 VSS.n40 VSS.t139 165.032
R3040 VSS.n39 VSS.t88 165.032
R3041 VSS.n38 VSS.t94 165.032
R3042 VSS.n37 VSS.t49 165.032
R3043 VSS.n36 VSS.t41 165.032
R3044 VSS.n35 VSS.t161 165.032
R3045 VSS.n34 VSS.t163 165.032
R3046 VSS.n33 VSS.t159 165.032
R3047 VSS.n32 VSS.t86 165.032
R3048 VSS.n400 VSS.t36 163.058
R3049 VSS.n402 VSS.t83 163.058
R3050 VSS.n404 VSS.t38 163.058
R3051 VSS.n406 VSS.t149 163.058
R3052 VSS.n408 VSS.t151 163.058
R3053 VSS.n397 VSS.t113 163.058
R3054 VSS.n411 VSS.t124 163.058
R3055 VSS.n394 VSS.t74 163.058
R3056 VSS.n392 VSS.t77 163.058
R3057 VSS.n390 VSS.t80 163.058
R3058 VSS.n388 VSS.t117 163.058
R3059 VSS.n386 VSS.t34 163.058
R3060 VSS.n413 VSS.t25 162.941
R3061 VSS.n413 VSS.t169 162.941
R3062 VSS.n400 VSS.t12 162.781
R3063 VSS.n402 VSS.t143 162.781
R3064 VSS.n404 VSS.t119 162.781
R3065 VSS.n406 VSS.t56 162.781
R3066 VSS.n408 VSS.t62 162.781
R3067 VSS.n394 VSS.t137 162.781
R3068 VSS.n392 VSS.t141 162.781
R3069 VSS.n390 VSS.t133 162.781
R3070 VSS.n388 VSS.t53 162.781
R3071 VSS.n386 VSS.t104 162.781
R3072 VSS.t25 VSS.n412 162.639
R3073 VSS.n396 VSS.t169 162.639
R3074 VSS.n1455 VSS.n1168 157.957
R3075 VSS.n283 VSS.n282 147.374
R3076 VSS.n290 VSS.n289 147.374
R3077 VSS.n291 VSS.n280 147.374
R3078 VSS.n298 VSS.n297 147.374
R3079 VSS.n299 VSS.n278 147.374
R3080 VSS.n306 VSS.n305 147.374
R3081 VSS.n307 VSS.n276 147.374
R3082 VSS.n314 VSS.n313 147.374
R3083 VSS.n315 VSS.n274 147.374
R3084 VSS.n322 VSS.n321 147.374
R3085 VSS.n323 VSS.n270 147.374
R3086 VSS.n484 VSS.n483 147.374
R3087 VSS.n485 VSS.n268 147.374
R3088 VSS.n492 VSS.n491 147.374
R3089 VSS.n493 VSS.n266 147.374
R3090 VSS.n500 VSS.n499 147.374
R3091 VSS.n501 VSS.n264 147.374
R3092 VSS.n508 VSS.n507 147.374
R3093 VSS.n509 VSS.n262 147.374
R3094 VSS.n2541 VSS.n2540 147.374
R3095 VSS.n2535 VSS.n122 147.374
R3096 VSS.n2532 VSS.n123 147.374
R3097 VSS.n2528 VSS.n124 147.374
R3098 VSS.n2524 VSS.n125 147.374
R3099 VSS.n2520 VSS.n126 147.374
R3100 VSS.n2516 VSS.n127 147.374
R3101 VSS.n2512 VSS.n128 147.374
R3102 VSS.n2508 VSS.n129 147.374
R3103 VSS.n2504 VSS.n130 147.374
R3104 VSS.n2495 VSS.n131 147.374
R3105 VSS.n2543 VSS.n120 147.374
R3106 VSS.n132 VSS.n119 147.374
R3107 VSS.n2462 VSS.n133 147.374
R3108 VSS.n2466 VSS.n134 147.374
R3109 VSS.n2470 VSS.n135 147.374
R3110 VSS.n2474 VSS.n136 147.374
R3111 VSS.n2478 VSS.n137 147.374
R3112 VSS.n2482 VSS.n138 147.374
R3113 VSS.n1782 VSS.n1735 147.374
R3114 VSS.n1778 VSS.n1734 147.374
R3115 VSS.n1774 VSS.n1733 147.374
R3116 VSS.n1770 VSS.n1732 147.374
R3117 VSS.n1766 VSS.n1731 147.374
R3118 VSS.n1762 VSS.n1730 147.374
R3119 VSS.n1758 VSS.n1729 147.374
R3120 VSS.n1754 VSS.n1728 147.374
R3121 VSS.n1750 VSS.n1727 147.374
R3122 VSS.n1746 VSS.n1726 147.374
R3123 VSS.n1742 VSS.n1725 147.374
R3124 VSS.n1862 VSS.n836 147.374
R3125 VSS.n1860 VSS.n839 147.374
R3126 VSS.n1856 VSS.n1855 147.374
R3127 VSS.n1849 VSS.n841 147.374
R3128 VSS.n1848 VSS.n1847 147.374
R3129 VSS.n1839 VSS.n843 147.374
R3130 VSS.n1838 VSS.n1837 147.374
R3131 VSS.n1831 VSS.n846 147.374
R3132 VSS.n1830 VSS.n1829 147.374
R3133 VSS.n1823 VSS.n848 147.374
R3134 VSS.n1822 VSS.n1821 147.374
R3135 VSS.n1288 VSS.n1287 147.374
R3136 VSS.n1285 VSS.n1284 147.374
R3137 VSS.n1280 VSS.n1241 147.374
R3138 VSS.n1278 VSS.n1277 147.374
R3139 VSS.n1273 VSS.n1244 147.374
R3140 VSS.n1271 VSS.n1270 147.374
R3141 VSS.n1266 VSS.n1247 147.374
R3142 VSS.n1264 VSS.n1263 147.374
R3143 VSS.n1259 VSS.n1250 147.374
R3144 VSS.n1257 VSS.n1256 147.374
R3145 VSS.n1251 VSS.n1235 147.374
R3146 VSS.n1590 VSS.n1589 147.374
R3147 VSS.n1584 VSS.n1081 147.374
R3148 VSS.n1581 VSS.n1082 147.374
R3149 VSS.n1577 VSS.n1083 147.374
R3150 VSS.n1573 VSS.n1084 147.374
R3151 VSS.n1569 VSS.n1085 147.374
R3152 VSS.n1565 VSS.n1086 147.374
R3153 VSS.n1561 VSS.n1087 147.374
R3154 VSS.n1557 VSS.n1088 147.374
R3155 VSS.n1553 VSS.n1089 147.374
R3156 VSS.n1549 VSS.n1090 147.374
R3157 VSS.n1132 VSS.n1120 147.374
R3158 VSS.n1136 VSS.n1121 147.374
R3159 VSS.n1140 VSS.n1122 147.374
R3160 VSS.n1144 VSS.n1123 147.374
R3161 VSS.n1148 VSS.n1124 147.374
R3162 VSS.n1152 VSS.n1125 147.374
R3163 VSS.n1156 VSS.n1126 147.374
R3164 VSS.n1160 VSS.n1127 147.374
R3165 VSS.n1163 VSS.n1128 147.374
R3166 VSS.n1462 VSS.n1461 147.374
R3167 VSS.n1457 VSS.n1167 147.374
R3168 VSS.n1450 VSS.n1171 147.374
R3169 VSS.n1448 VSS.n1447 147.374
R3170 VSS.n1443 VSS.n1174 147.374
R3171 VSS.n1441 VSS.n1440 147.374
R3172 VSS.n1436 VSS.n1177 147.374
R3173 VSS.n1434 VSS.n1433 147.374
R3174 VSS.n1429 VSS.n1180 147.374
R3175 VSS.n1427 VSS.n1426 147.374
R3176 VSS.n1422 VSS.n1183 147.374
R3177 VSS.n1420 VSS.n1419 147.374
R3178 VSS.n1415 VSS.n1186 147.374
R3179 VSS.n1408 VSS.n1189 147.374
R3180 VSS.n1406 VSS.n1405 147.374
R3181 VSS.n1401 VSS.n1192 147.374
R3182 VSS.n1399 VSS.n1398 147.374
R3183 VSS.n1394 VSS.n1195 147.374
R3184 VSS.n1392 VSS.n1391 147.374
R3185 VSS.n1387 VSS.n1198 147.374
R3186 VSS.n1385 VSS.n1384 147.374
R3187 VSS.n1380 VSS.n1201 147.374
R3188 VSS.n1378 VSS.n1377 147.374
R3189 VSS.n1373 VSS.n1204 147.374
R3190 VSS.n1366 VSS.n1207 147.374
R3191 VSS.n1364 VSS.n1363 147.374
R3192 VSS.n1359 VSS.n1210 147.374
R3193 VSS.n1357 VSS.n1356 147.374
R3194 VSS.n1352 VSS.n1213 147.374
R3195 VSS.n1350 VSS.n1349 147.374
R3196 VSS.n1345 VSS.n1216 147.374
R3197 VSS.n1343 VSS.n1342 147.374
R3198 VSS.n1338 VSS.n1219 147.374
R3199 VSS.n1336 VSS.n1335 147.374
R3200 VSS.n1331 VSS.n1222 147.374
R3201 VSS.n2064 VSS.n768 147.374
R3202 VSS.n2059 VSS.n770 147.374
R3203 VSS.n2056 VSS.n771 147.374
R3204 VSS.n2052 VSS.n772 147.374
R3205 VSS.n2048 VSS.n773 147.374
R3206 VSS.n2044 VSS.n774 147.374
R3207 VSS.n2040 VSS.n775 147.374
R3208 VSS.n2036 VSS.n776 147.374
R3209 VSS.n2032 VSS.n777 147.374
R3210 VSS.n2026 VSS.n2025 147.374
R3211 VSS.n822 VSS.n783 147.374
R3212 VSS.n2018 VSS.n784 147.374
R3213 VSS.n2014 VSS.n785 147.374
R3214 VSS.n2010 VSS.n786 147.374
R3215 VSS.n2006 VSS.n787 147.374
R3216 VSS.n2002 VSS.n788 147.374
R3217 VSS.n1998 VSS.n789 147.374
R3218 VSS.n1994 VSS.n790 147.374
R3219 VSS.n1990 VSS.n791 147.374
R3220 VSS.n1986 VSS.n792 147.374
R3221 VSS.n1982 VSS.n793 147.374
R3222 VSS.n1978 VSS.n794 147.374
R3223 VSS.n1974 VSS.n795 147.374
R3224 VSS.n1970 VSS.n796 147.374
R3225 VSS.n1966 VSS.n797 147.374
R3226 VSS.n1962 VSS.n798 147.374
R3227 VSS.n1958 VSS.n799 147.374
R3228 VSS.n1954 VSS.n800 147.374
R3229 VSS.n1950 VSS.n801 147.374
R3230 VSS.n1946 VSS.n802 147.374
R3231 VSS.n1942 VSS.n803 147.374
R3232 VSS.n1938 VSS.n804 147.374
R3233 VSS.n1934 VSS.n805 147.374
R3234 VSS.n1930 VSS.n806 147.374
R3235 VSS.n1926 VSS.n807 147.374
R3236 VSS.n1922 VSS.n808 147.374
R3237 VSS.n1918 VSS.n809 147.374
R3238 VSS.n1914 VSS.n810 147.374
R3239 VSS.n1910 VSS.n811 147.374
R3240 VSS.n1906 VSS.n812 147.374
R3241 VSS.n1902 VSS.n813 147.374
R3242 VSS.n1898 VSS.n814 147.374
R3243 VSS.n1894 VSS.n815 147.374
R3244 VSS.n1890 VSS.n816 147.374
R3245 VSS.n1886 VSS.n817 147.374
R3246 VSS.n2112 VSS.n642 147.374
R3247 VSS.n2110 VSS.n644 147.374
R3248 VSS.n2282 VSS.n529 147.374
R3249 VSS.n2278 VSS.n528 147.374
R3250 VSS.n2281 VSS.n528 147.374
R3251 VSS.n531 VSS.n529 147.374
R3252 VSS.n2113 VSS.n2112 147.374
R3253 VSS.n644 VSS.n640 147.374
R3254 VSS.n2064 VSS.n2063 147.374
R3255 VSS.n2057 VSS.n770 147.374
R3256 VSS.n2053 VSS.n771 147.374
R3257 VSS.n2049 VSS.n772 147.374
R3258 VSS.n2045 VSS.n773 147.374
R3259 VSS.n2041 VSS.n774 147.374
R3260 VSS.n2037 VSS.n775 147.374
R3261 VSS.n2033 VSS.n776 147.374
R3262 VSS.n2029 VSS.n777 147.374
R3263 VSS.n1462 VSS.n1129 147.374
R3264 VSS.n1161 VSS.n1128 147.374
R3265 VSS.n1157 VSS.n1127 147.374
R3266 VSS.n1153 VSS.n1126 147.374
R3267 VSS.n1149 VSS.n1125 147.374
R3268 VSS.n1145 VSS.n1124 147.374
R3269 VSS.n1141 VSS.n1123 147.374
R3270 VSS.n1137 VSS.n1122 147.374
R3271 VSS.n1133 VSS.n1121 147.374
R3272 VSS.n1120 VSS.n1119 147.374
R3273 VSS.n1590 VSS.n1092 147.374
R3274 VSS.n1582 VSS.n1081 147.374
R3275 VSS.n1578 VSS.n1082 147.374
R3276 VSS.n1574 VSS.n1083 147.374
R3277 VSS.n1570 VSS.n1084 147.374
R3278 VSS.n1566 VSS.n1085 147.374
R3279 VSS.n1562 VSS.n1086 147.374
R3280 VSS.n1558 VSS.n1087 147.374
R3281 VSS.n1554 VSS.n1088 147.374
R3282 VSS.n1550 VSS.n1089 147.374
R3283 VSS.n1546 VSS.n1090 147.374
R3284 VSS.n1252 VSS.n1251 147.374
R3285 VSS.n1258 VSS.n1257 147.374
R3286 VSS.n1250 VSS.n1248 147.374
R3287 VSS.n1265 VSS.n1264 147.374
R3288 VSS.n1247 VSS.n1245 147.374
R3289 VSS.n1272 VSS.n1271 147.374
R3290 VSS.n1244 VSS.n1242 147.374
R3291 VSS.n1279 VSS.n1278 147.374
R3292 VSS.n1241 VSS.n1239 147.374
R3293 VSS.n1286 VSS.n1285 147.374
R3294 VSS.n1289 VSS.n1288 147.374
R3295 VSS.n1863 VSS.n1862 147.374
R3296 VSS.n1857 VSS.n839 147.374
R3297 VSS.n1855 VSS.n1854 147.374
R3298 VSS.n1850 VSS.n1849 147.374
R3299 VSS.n1847 VSS.n1846 147.374
R3300 VSS.n1840 VSS.n1839 147.374
R3301 VSS.n1837 VSS.n1836 147.374
R3302 VSS.n1832 VSS.n1831 147.374
R3303 VSS.n1829 VSS.n1828 147.374
R3304 VSS.n1824 VSS.n1823 147.374
R3305 VSS.n1821 VSS.n1820 147.374
R3306 VSS.n1745 VSS.n1725 147.374
R3307 VSS.n1749 VSS.n1726 147.374
R3308 VSS.n1753 VSS.n1727 147.374
R3309 VSS.n1757 VSS.n1728 147.374
R3310 VSS.n1761 VSS.n1729 147.374
R3311 VSS.n1765 VSS.n1730 147.374
R3312 VSS.n1769 VSS.n1731 147.374
R3313 VSS.n1773 VSS.n1732 147.374
R3314 VSS.n1777 VSS.n1733 147.374
R3315 VSS.n1781 VSS.n1734 147.374
R3316 VSS.n1736 VSS.n1735 147.374
R3317 VSS.n2541 VSS.n141 147.374
R3318 VSS.n2533 VSS.n122 147.374
R3319 VSS.n2529 VSS.n123 147.374
R3320 VSS.n2525 VSS.n124 147.374
R3321 VSS.n2521 VSS.n125 147.374
R3322 VSS.n2517 VSS.n126 147.374
R3323 VSS.n2513 VSS.n127 147.374
R3324 VSS.n2509 VSS.n128 147.374
R3325 VSS.n2505 VSS.n129 147.374
R3326 VSS.n2494 VSS.n130 147.374
R3327 VSS.n2498 VSS.n131 147.374
R3328 VSS.n2544 VSS.n2543 147.374
R3329 VSS.n2461 VSS.n132 147.374
R3330 VSS.n2465 VSS.n133 147.374
R3331 VSS.n2469 VSS.n134 147.374
R3332 VSS.n2473 VSS.n135 147.374
R3333 VSS.n2477 VSS.n136 147.374
R3334 VSS.n2481 VSS.n137 147.374
R3335 VSS.n2484 VSS.n138 147.374
R3336 VSS.n510 VSS.n509 147.374
R3337 VSS.n507 VSS.n506 147.374
R3338 VSS.n502 VSS.n501 147.374
R3339 VSS.n499 VSS.n498 147.374
R3340 VSS.n494 VSS.n493 147.374
R3341 VSS.n491 VSS.n490 147.374
R3342 VSS.n486 VSS.n485 147.374
R3343 VSS.n483 VSS.n482 147.374
R3344 VSS.n324 VSS.n323 147.374
R3345 VSS.n321 VSS.n320 147.374
R3346 VSS.n316 VSS.n315 147.374
R3347 VSS.n313 VSS.n312 147.374
R3348 VSS.n308 VSS.n307 147.374
R3349 VSS.n305 VSS.n304 147.374
R3350 VSS.n300 VSS.n299 147.374
R3351 VSS.n297 VSS.n296 147.374
R3352 VSS.n292 VSS.n291 147.374
R3353 VSS.n289 VSS.n288 147.374
R3354 VSS.n284 VSS.n283 147.374
R3355 VSS.n2025 VSS.n781 147.374
R3356 VSS.n2019 VSS.n783 147.374
R3357 VSS.n2015 VSS.n784 147.374
R3358 VSS.n2011 VSS.n785 147.374
R3359 VSS.n2007 VSS.n786 147.374
R3360 VSS.n2003 VSS.n787 147.374
R3361 VSS.n1999 VSS.n788 147.374
R3362 VSS.n1995 VSS.n789 147.374
R3363 VSS.n1991 VSS.n790 147.374
R3364 VSS.n1987 VSS.n791 147.374
R3365 VSS.n1983 VSS.n792 147.374
R3366 VSS.n1979 VSS.n793 147.374
R3367 VSS.n1975 VSS.n794 147.374
R3368 VSS.n1971 VSS.n795 147.374
R3369 VSS.n1967 VSS.n796 147.374
R3370 VSS.n1963 VSS.n797 147.374
R3371 VSS.n1959 VSS.n798 147.374
R3372 VSS.n1955 VSS.n799 147.374
R3373 VSS.n1951 VSS.n800 147.374
R3374 VSS.n1947 VSS.n801 147.374
R3375 VSS.n1943 VSS.n802 147.374
R3376 VSS.n1939 VSS.n803 147.374
R3377 VSS.n1935 VSS.n804 147.374
R3378 VSS.n1931 VSS.n805 147.374
R3379 VSS.n1927 VSS.n806 147.374
R3380 VSS.n1923 VSS.n807 147.374
R3381 VSS.n1919 VSS.n808 147.374
R3382 VSS.n1915 VSS.n809 147.374
R3383 VSS.n1911 VSS.n810 147.374
R3384 VSS.n1907 VSS.n811 147.374
R3385 VSS.n1903 VSS.n812 147.374
R3386 VSS.n1899 VSS.n813 147.374
R3387 VSS.n1895 VSS.n814 147.374
R3388 VSS.n1891 VSS.n815 147.374
R3389 VSS.n1887 VSS.n816 147.374
R3390 VSS.n1883 VSS.n817 147.374
R3391 VSS.n1222 VSS.n1220 147.374
R3392 VSS.n1337 VSS.n1336 147.374
R3393 VSS.n1219 VSS.n1217 147.374
R3394 VSS.n1344 VSS.n1343 147.374
R3395 VSS.n1216 VSS.n1214 147.374
R3396 VSS.n1351 VSS.n1350 147.374
R3397 VSS.n1213 VSS.n1211 147.374
R3398 VSS.n1358 VSS.n1357 147.374
R3399 VSS.n1210 VSS.n1208 147.374
R3400 VSS.n1365 VSS.n1364 147.374
R3401 VSS.n1207 VSS.n1205 147.374
R3402 VSS.n1204 VSS.n1202 147.374
R3403 VSS.n1379 VSS.n1378 147.374
R3404 VSS.n1201 VSS.n1199 147.374
R3405 VSS.n1386 VSS.n1385 147.374
R3406 VSS.n1198 VSS.n1196 147.374
R3407 VSS.n1393 VSS.n1392 147.374
R3408 VSS.n1195 VSS.n1193 147.374
R3409 VSS.n1400 VSS.n1399 147.374
R3410 VSS.n1192 VSS.n1190 147.374
R3411 VSS.n1407 VSS.n1406 147.374
R3412 VSS.n1189 VSS.n1187 147.374
R3413 VSS.n1186 VSS.n1184 147.374
R3414 VSS.n1421 VSS.n1420 147.374
R3415 VSS.n1183 VSS.n1181 147.374
R3416 VSS.n1428 VSS.n1427 147.374
R3417 VSS.n1180 VSS.n1178 147.374
R3418 VSS.n1435 VSS.n1434 147.374
R3419 VSS.n1177 VSS.n1175 147.374
R3420 VSS.n1442 VSS.n1441 147.374
R3421 VSS.n1174 VSS.n1172 147.374
R3422 VSS.n1449 VSS.n1448 147.374
R3423 VSS.n1171 VSS.n1169 147.374
R3424 VSS.n1167 VSS.n1130 147.374
R3425 VSS.n1716 VSS.n1715 147.374
R3426 VSS.n1710 VSS.n869 147.374
R3427 VSS.n1707 VSS.n870 147.374
R3428 VSS.n1703 VSS.n871 147.374
R3429 VSS.n1699 VSS.n872 147.374
R3430 VSS.n1695 VSS.n873 147.374
R3431 VSS.n1691 VSS.n874 147.374
R3432 VSS.n1687 VSS.n875 147.374
R3433 VSS.n1683 VSS.n876 147.374
R3434 VSS.n1679 VSS.n877 147.374
R3435 VSS.n1675 VSS.n878 147.374
R3436 VSS.n1602 VSS.n1023 147.374
R3437 VSS.n1028 VSS.n1027 147.374
R3438 VSS.n1040 VSS.n1029 147.374
R3439 VSS.n1044 VSS.n1030 147.374
R3440 VSS.n1048 VSS.n1031 147.374
R3441 VSS.n1052 VSS.n1032 147.374
R3442 VSS.n1056 VSS.n1033 147.374
R3443 VSS.n1060 VSS.n1034 147.374
R3444 VSS.n1064 VSS.n1035 147.374
R3445 VSS.n1068 VSS.n1036 147.374
R3446 VSS.n1075 VSS.n1037 147.374
R3447 VSS.n1075 VSS.n1074 147.374
R3448 VSS.n1070 VSS.n1036 147.374
R3449 VSS.n1067 VSS.n1035 147.374
R3450 VSS.n1063 VSS.n1034 147.374
R3451 VSS.n1059 VSS.n1033 147.374
R3452 VSS.n1055 VSS.n1032 147.374
R3453 VSS.n1051 VSS.n1031 147.374
R3454 VSS.n1047 VSS.n1030 147.374
R3455 VSS.n1043 VSS.n1029 147.374
R3456 VSS.n1039 VSS.n1028 147.374
R3457 VSS.n1603 VSS.n1602 147.374
R3458 VSS.n1716 VSS.n880 147.374
R3459 VSS.n1708 VSS.n869 147.374
R3460 VSS.n1704 VSS.n870 147.374
R3461 VSS.n1700 VSS.n871 147.374
R3462 VSS.n1696 VSS.n872 147.374
R3463 VSS.n1692 VSS.n873 147.374
R3464 VSS.n1688 VSS.n874 147.374
R3465 VSS.n1684 VSS.n875 147.374
R3466 VSS.n1680 VSS.n876 147.374
R3467 VSS.n1676 VSS.n877 147.374
R3468 VSS.n1672 VSS.n878 147.374
R3469 VSS.n111 VSS.n87 140.69
R3470 VSS.n104 VSS.n87 140.69
R3471 VSS.n58 VSS.n57 140.69
R3472 VSS.n58 VSS.n49 140.69
R3473 VSS.n979 VSS.n973 140.69
R3474 VSS.n980 VSS.n979 140.69
R3475 VSS.n980 VSS.n969 140.69
R3476 VSS.n987 VSS.n969 140.69
R3477 VSS.n988 VSS.n987 140.69
R3478 VSS.n988 VSS.n965 140.69
R3479 VSS.n995 VSS.n965 140.69
R3480 VSS.n954 VSS.n921 140.69
R3481 VSS.n947 VSS.n921 140.69
R3482 VSS.n947 VSS.n946 140.69
R3483 VSS.n946 VSS.n925 140.69
R3484 VSS.n939 VSS.n925 140.69
R3485 VSS.n939 VSS.n938 140.69
R3486 VSS.n938 VSS.n929 140.69
R3487 VSS.n730 VSS.n729 140.69
R3488 VSS.n729 VSS.n703 140.69
R3489 VSS.n722 VSS.n703 140.69
R3490 VSS.n722 VSS.n721 140.69
R3491 VSS.n721 VSS.n707 140.69
R3492 VSS.n714 VSS.n707 140.69
R3493 VSS.n714 VSS.n713 140.69
R3494 VSS.n670 VSS.n664 140.69
R3495 VSS.n677 VSS.n664 140.69
R3496 VSS.n678 VSS.n677 140.69
R3497 VSS.n678 VSS.n660 140.69
R3498 VSS.n686 VSS.n660 140.69
R3499 VSS.n687 VSS.n686 140.69
R3500 VSS.n687 VSS.n657 140.69
R3501 VSS.n13 VSS.t90 130.75
R3502 VSS.n1465 VSS.n1463 120.079
R3503 VSS.n2066 VSS.n2065 120.079
R3504 VSS.n2118 VSS.n637 109.478
R3505 VSS.n2124 VSS.n637 109.478
R3506 VSS.n2124 VSS.n633 109.478
R3507 VSS.n2130 VSS.n633 109.478
R3508 VSS.n2130 VSS.n629 109.478
R3509 VSS.n2136 VSS.n629 109.478
R3510 VSS.n2136 VSS.n625 109.478
R3511 VSS.n2142 VSS.n625 109.478
R3512 VSS.n2142 VSS.n621 109.478
R3513 VSS.n2148 VSS.n621 109.478
R3514 VSS.n2148 VSS.n616 109.478
R3515 VSS.n2154 VSS.n616 109.478
R3516 VSS.n2160 VSS.n612 109.478
R3517 VSS.n2160 VSS.n608 109.478
R3518 VSS.n2166 VSS.n608 109.478
R3519 VSS.n2166 VSS.n604 109.478
R3520 VSS.n2172 VSS.n604 109.478
R3521 VSS.n2172 VSS.n600 109.478
R3522 VSS.n2178 VSS.n600 109.478
R3523 VSS.n2178 VSS.n596 109.478
R3524 VSS.n2184 VSS.n596 109.478
R3525 VSS.n2184 VSS.n592 109.478
R3526 VSS.n2190 VSS.n592 109.478
R3527 VSS.n2190 VSS.n588 109.478
R3528 VSS.n2196 VSS.n588 109.478
R3529 VSS.n2202 VSS.n584 109.478
R3530 VSS.n2202 VSS.n580 109.478
R3531 VSS.n2208 VSS.n580 109.478
R3532 VSS.n2208 VSS.n576 109.478
R3533 VSS.n2214 VSS.n576 109.478
R3534 VSS.n2214 VSS.n572 109.478
R3535 VSS.n2220 VSS.n572 109.478
R3536 VSS.n2220 VSS.n568 109.478
R3537 VSS.n2226 VSS.n568 109.478
R3538 VSS.n2226 VSS.n564 109.478
R3539 VSS.n2232 VSS.n564 109.478
R3540 VSS.n2232 VSS.n560 109.478
R3541 VSS.n2238 VSS.n560 109.478
R3542 VSS.n2238 VSS.n556 109.478
R3543 VSS.n2244 VSS.n556 109.478
R3544 VSS.n2244 VSS.n552 109.478
R3545 VSS.n2250 VSS.n552 109.478
R3546 VSS.n2250 VSS.n548 109.478
R3547 VSS.n2256 VSS.n548 109.478
R3548 VSS.n2256 VSS.n544 109.478
R3549 VSS.n2262 VSS.n544 109.478
R3550 VSS.n2262 VSS.n540 109.478
R3551 VSS.n2269 VSS.n540 109.478
R3552 VSS.n2269 VSS.n536 109.478
R3553 VSS.n2275 VSS.n536 109.478
R3554 VSS.n2275 VSS.n527 109.478
R3555 VSS.n13 VSS.t93 91.3557
R3556 VSS.n362 VSS.t61 90.6265
R3557 VSS.n346 VSS.t33 90.6265
R3558 VSS.n461 VSS.t99 90.6265
R3559 VSS.n444 VSS.t67 90.6265
R3560 VSS.n428 VSS.n333 86.5152
R3561 VSS.n30 VSS.n29 86.5152
R3562 VSS.n2116 VSS.n2115 85.8358
R3563 VSS.n2285 VSS.n532 85.8358
R3564 VSS.n2279 VSS.n533 85.8358
R3565 VSS.n1785 VSS.n855 82.4476
R3566 VSS.n1866 VSS.n1865 82.4476
R3567 VSS.n1743 VSS.n1739 82.4476
R3568 VSS.n1819 VSS.n1818 82.4476
R3569 VSS.n1292 VSS.n1291 82.4476
R3570 VSS.n1588 VSS.n1094 82.4476
R3571 VSS.n1253 VSS.n1234 82.4476
R3572 VSS.n1547 VSS.n1095 82.4476
R3573 VSS.n1607 VSS.n1605 82.4476
R3574 VSS.n1611 VSS.n1019 82.4476
R3575 VSS.n1714 VSS.n882 82.4476
R3576 VSS.n1673 VSS.n883 82.4476
R3577 VSS.n362 VSS.t59 81.8918
R3578 VSS.n361 VSS.t157 81.8918
R3579 VSS.n346 VSS.t30 81.8918
R3580 VSS.n465 VSS.t96 81.8918
R3581 VSS.n461 VSS.t98 81.8918
R3582 VSS.n444 VSS.t65 81.8918
R3583 VSS.n89 VSS.t71 81.8918
R3584 VSS.n102 VSS.t126 81.8918
R3585 VSS.n48 VSS.t155 81.8918
R3586 VSS.n65 VSS.t153 81.8918
R3587 VSS.n617 VSS.n612 80.4981
R3588 VSS.n517 VSS.n259 76.8005
R3589 VSS.n2539 VSS.n2492 76.8005
R3590 VSS.n513 VSS.n512 76.8005
R3591 VSS.n2486 VSS.n2485 76.8005
R3592 VSS.n1467 VSS.n1118 76.8005
R3593 VSS.n2068 VSS.n767 76.8005
R3594 VSS.n1332 VSS.n1221 76.8005
R3595 VSS.n1882 VSS.n1881 76.8005
R3596 VSS.n1465 VSS.n1464 72.905
R3597 VSS.n1472 VSS.n1471 72.905
R3598 VSS.n1473 VSS.n1472 72.905
R3599 VSS.n1473 VSS.n1111 72.905
R3600 VSS.n1518 VSS.n1112 72.905
R3601 VSS.n1512 VSS.n1112 72.905
R3602 VSS.n1512 VSS.n1098 72.905
R3603 VSS.n1503 VSS.n1099 72.905
R3604 VSS.n1505 VSS.n1503 72.905
R3605 VSS.n1505 VSS.n1504 72.905
R3606 VSS.n1500 VSS.n1499 72.905
R3607 VSS.n1499 VSS.n1498 72.905
R3608 VSS.n1489 VSS.n1017 72.905
R3609 VSS.n1489 VSS.n1488 72.905
R3610 VSS.n2098 VSS.n752 72.905
R3611 VSS.n2098 VSS.n2097 72.905
R3612 VSS.n2097 VSS.n2096 72.905
R3613 VSS.n2090 VSS.n757 72.905
R3614 VSS.n2090 VSS.n2089 72.905
R3615 VSS.n2089 VSS.n2088 72.905
R3616 VSS.n2082 VSS.n761 72.905
R3617 VSS.n2082 VSS.n2081 72.905
R3618 VSS.n2081 VSS.n2080 72.905
R3619 VSS.n2074 VSS.n765 72.905
R3620 VSS.n2074 VSS.n2073 72.905
R3621 VSS.n2073 VSS.n2072 72.905
R3622 VSS.n2066 VSS.n769 72.905
R3623 VSS.n104 VSS.t128 70.3453
R3624 VSS.t156 VSS.n49 70.3453
R3625 VSS.t24 VSS.n973 70.3453
R3626 VSS.t29 VSS.n954 70.3453
R3627 VSS.n713 VSS.t123 70.3453
R3628 VSS.t19 VSS.n657 70.3453
R3629 VSS.n1464 VSS.t9 67.5444
R3630 VSS.n769 VSS.t8 67.5444
R3631 VSS.n1868 VSS.n835 66.162
R3632 VSS.t111 VSS.n1017 65.4001
R3633 VSS.n1488 VSS.t7 65.4001
R3634 VSS.n1453 VSS.n1166 64.7534
R3635 VSS.n2022 VSS.n2021 64.7534
R3636 VSS.n2120 VSS.n639 62.1181
R3637 VSS.n1168 VSS.n139 61.9943
R3638 VSS.n1498 VSS.n1015 57.8952
R3639 VSS.n2196 VSS.t175 54.7389
R3640 VSS.t175 VSS.n584 54.7389
R3641 VSS.n515 VSS.n261 54.18
R3642 VSS.n2542 VSS.n121 54.18
R3643 VSS.t1 VSS.n1111 52.5346
R3644 VSS.n765 VSS.t5 52.5346
R3645 VSS.n1500 VSS.t0 50.3904
R3646 VSS.n2096 VSS.t45 50.3904
R3647 VSS.n1411 VSS.n1185 39.1534
R3648 VSS.n1369 VSS.n1203 39.1534
R3649 VSS.n1976 VSS.n1973 39.1534
R3650 VSS.n1928 VSS.n1925 39.1534
R3651 VSS.t2 VSS.n1098 37.5249
R3652 VSS.n761 VSS.t4 37.5249
R3653 VSS.n515 VSS.n257 35.4256
R3654 VSS.n521 VSS.n257 35.4256
R3655 VSS.n2290 VSS.n253 35.4256
R3656 VSS.n2296 VSS.n246 35.4256
R3657 VSS.n2303 VSS.n246 35.4256
R3658 VSS.n2303 VSS.n2302 35.4256
R3659 VSS.n2309 VSS.n239 35.4256
R3660 VSS.n2316 VSS.n239 35.4256
R3661 VSS.n2316 VSS.n2315 35.4256
R3662 VSS.n2322 VSS.n232 35.4256
R3663 VSS.n2329 VSS.n232 35.4256
R3664 VSS.n2329 VSS.n2328 35.4256
R3665 VSS.n2335 VSS.n225 35.4256
R3666 VSS.n2342 VSS.n225 35.4256
R3667 VSS.n2342 VSS.n2341 35.4256
R3668 VSS.n2348 VSS.n218 35.4256
R3669 VSS.n2354 VSS.n218 35.4256
R3670 VSS.n2360 VSS.n214 35.4256
R3671 VSS.n2360 VSS.n210 35.4256
R3672 VSS.n2366 VSS.n210 35.4256
R3673 VSS.n2372 VSS.n206 35.4256
R3674 VSS.n2372 VSS.n202 35.4256
R3675 VSS.n2378 VSS.n202 35.4256
R3676 VSS.n2384 VSS.n198 35.4256
R3677 VSS.n2384 VSS.n194 35.4256
R3678 VSS.n2390 VSS.n194 35.4256
R3679 VSS.n2396 VSS.n189 35.4256
R3680 VSS.n2396 VSS.n190 35.4256
R3681 VSS.n2402 VSS.n181 35.4256
R3682 VSS.n2408 VSS.n181 35.4256
R3683 VSS.n2408 VSS.n182 35.4256
R3684 VSS.n2414 VSS.n173 35.4256
R3685 VSS.n2420 VSS.n173 35.4256
R3686 VSS.n2420 VSS.n174 35.4256
R3687 VSS.n2426 VSS.n165 35.4256
R3688 VSS.n2432 VSS.n165 35.4256
R3689 VSS.n2432 VSS.n166 35.4256
R3690 VSS.n2438 VSS.n157 35.4256
R3691 VSS.n2444 VSS.n157 35.4256
R3692 VSS.n2444 VSS.n158 35.4256
R3693 VSS.n2450 VSS.n150 35.4256
R3694 VSS.n2456 VSS.n150 35.4256
R3695 VSS.n2489 VSS.n145 35.4256
R3696 VSS.n2489 VSS.n121 35.4256
R3697 VSS.n1294 VSS.n1224 35.4256
R3698 VSS.n1543 VSS.n1080 35.4256
R3699 VSS.n1593 VSS.n1592 35.4256
R3700 VSS.n1600 VSS.n1021 35.4256
R3701 VSS.n1718 VSS.n868 35.4256
R3702 VSS.n1724 VSS.n864 35.4256
R3703 VSS.n1789 VSS.n1788 35.4256
R3704 VSS.n2024 VSS.n782 35.4256
R3705 VSS.n2024 VSS.n820 35.4256
R3706 VSS.n1870 VSS.n820 35.4256
R3707 VSS.n1869 VSS.n1868 35.4256
R3708 VSS.t2 VSS.n1099 35.3806
R3709 VSS.n2088 VSS.t4 35.3806
R3710 VSS.n2348 VSS.t78 34.9046
R3711 VSS.n190 VSS.t57 34.9046
R3712 VSS.t66 VSS.n253 33.8627
R3713 VSS.n2456 VSS.t31 33.8627
R3714 VSS.n353 VSS.n352 32.8962
R3715 VSS.n451 VSS.n450 32.8962
R3716 VSS.n2289 VSS.n2288 30.7369
R3717 VSS.n28 VSS.n12 30.3012
R3718 VSS.n2288 VSS.t69 29.695
R3719 VSS.n2450 VSS.t72 29.695
R3720 VSS.n2154 VSS.n617 28.9796
R3721 VSS.n2354 VSS.t75 28.6531
R3722 VSS.t63 VSS.n189 28.6531
R3723 VSS.n105 VSS.n103 28.3989
R3724 VSS.n62 VSS.n61 28.3989
R3725 VSS.n377 VSS.n376 27.9576
R3726 VSS.n381 VSS.n380 27.9576
R3727 VSS.n329 VSS.n328 27.9576
R3728 VSS.n432 VSS.n431 27.9576
R3729 VSS.n436 VSS.n435 27.9576
R3730 VSS.n375 VSS.n374 27.7293
R3731 VSS.n379 VSS.n378 27.7293
R3732 VSS.n383 VSS.n382 27.7293
R3733 VSS.n430 VSS.n429 27.7293
R3734 VSS.n434 VSS.n433 27.7293
R3735 VSS.n438 VSS.n437 27.7293
R3736 VSS.n83 VSS.n82 27.7293
R3737 VSS.n81 VSS.n80 27.7293
R3738 VSS.n79 VSS.n78 27.7293
R3739 VSS.n77 VSS.n76 27.7293
R3740 VSS.n75 VSS.n74 27.7293
R3741 VSS.n2335 VSS.t81 27.6112
R3742 VSS.n182 VSS.t39 27.6112
R3743 VSS.n1787 VSS.n1724 27.6112
R3744 VSS.n369 VSS.n340 27.5286
R3745 VSS.n370 VSS.n338 27.5286
R3746 VSS.n473 VSS.n456 27.5286
R3747 VSS.n472 VSS.n458 27.5286
R3748 VSS.n99 VSS.n90 27.5286
R3749 VSS.n70 VSS.n47 27.5286
R3750 VSS.n997 VSS.n996 25.6009
R3751 VSS.n932 VSS.n931 25.6009
R3752 VSS.n734 VSS.n700 25.6009
R3753 VSS.n669 VSS.n668 25.6009
R3754 VSS.n518 VSS.n517 25.6005
R3755 VSS.n519 VSS.n518 25.6005
R3756 VSS.n519 VSS.n251 25.6005
R3757 VSS.n2292 VSS.n251 25.6005
R3758 VSS.n2293 VSS.n2292 25.6005
R3759 VSS.n2294 VSS.n2293 25.6005
R3760 VSS.n2294 VSS.n244 25.6005
R3761 VSS.n2305 VSS.n244 25.6005
R3762 VSS.n2306 VSS.n2305 25.6005
R3763 VSS.n2307 VSS.n2306 25.6005
R3764 VSS.n2307 VSS.n237 25.6005
R3765 VSS.n2318 VSS.n237 25.6005
R3766 VSS.n2319 VSS.n2318 25.6005
R3767 VSS.n2320 VSS.n2319 25.6005
R3768 VSS.n2320 VSS.n230 25.6005
R3769 VSS.n2331 VSS.n230 25.6005
R3770 VSS.n2332 VSS.n2331 25.6005
R3771 VSS.n2333 VSS.n2332 25.6005
R3772 VSS.n2333 VSS.n223 25.6005
R3773 VSS.n2344 VSS.n223 25.6005
R3774 VSS.n2345 VSS.n2344 25.6005
R3775 VSS.n2346 VSS.n2345 25.6005
R3776 VSS.n2346 VSS.n216 25.6005
R3777 VSS.n2356 VSS.n216 25.6005
R3778 VSS.n2357 VSS.n2356 25.6005
R3779 VSS.n2358 VSS.n2357 25.6005
R3780 VSS.n2358 VSS.n208 25.6005
R3781 VSS.n2368 VSS.n208 25.6005
R3782 VSS.n2369 VSS.n2368 25.6005
R3783 VSS.n2370 VSS.n2369 25.6005
R3784 VSS.n2370 VSS.n200 25.6005
R3785 VSS.n2380 VSS.n200 25.6005
R3786 VSS.n2381 VSS.n2380 25.6005
R3787 VSS.n2382 VSS.n2381 25.6005
R3788 VSS.n2382 VSS.n192 25.6005
R3789 VSS.n2392 VSS.n192 25.6005
R3790 VSS.n2393 VSS.n2392 25.6005
R3791 VSS.n2394 VSS.n2393 25.6005
R3792 VSS.n2394 VSS.n184 25.6005
R3793 VSS.n2404 VSS.n184 25.6005
R3794 VSS.n2405 VSS.n2404 25.6005
R3795 VSS.n2406 VSS.n2405 25.6005
R3796 VSS.n2406 VSS.n176 25.6005
R3797 VSS.n2416 VSS.n176 25.6005
R3798 VSS.n2417 VSS.n2416 25.6005
R3799 VSS.n2418 VSS.n2417 25.6005
R3800 VSS.n2418 VSS.n168 25.6005
R3801 VSS.n2428 VSS.n168 25.6005
R3802 VSS.n2429 VSS.n2428 25.6005
R3803 VSS.n2430 VSS.n2429 25.6005
R3804 VSS.n2430 VSS.n160 25.6005
R3805 VSS.n2440 VSS.n160 25.6005
R3806 VSS.n2441 VSS.n2440 25.6005
R3807 VSS.n2442 VSS.n2441 25.6005
R3808 VSS.n2442 VSS.n152 25.6005
R3809 VSS.n2452 VSS.n152 25.6005
R3810 VSS.n2453 VSS.n2452 25.6005
R3811 VSS.n2454 VSS.n2453 25.6005
R3812 VSS.n2454 VSS.n143 25.6005
R3813 VSS.n2491 VSS.n143 25.6005
R3814 VSS.n2492 VSS.n2491 25.6005
R3815 VSS.n285 VSS.n259 25.6005
R3816 VSS.n286 VSS.n285 25.6005
R3817 VSS.n287 VSS.n286 25.6005
R3818 VSS.n287 VSS.n281 25.6005
R3819 VSS.n293 VSS.n281 25.6005
R3820 VSS.n294 VSS.n293 25.6005
R3821 VSS.n295 VSS.n294 25.6005
R3822 VSS.n295 VSS.n279 25.6005
R3823 VSS.n301 VSS.n279 25.6005
R3824 VSS.n302 VSS.n301 25.6005
R3825 VSS.n303 VSS.n302 25.6005
R3826 VSS.n303 VSS.n277 25.6005
R3827 VSS.n309 VSS.n277 25.6005
R3828 VSS.n310 VSS.n309 25.6005
R3829 VSS.n311 VSS.n310 25.6005
R3830 VSS.n311 VSS.n275 25.6005
R3831 VSS.n317 VSS.n275 25.6005
R3832 VSS.n318 VSS.n317 25.6005
R3833 VSS.n319 VSS.n318 25.6005
R3834 VSS.n325 VSS.n273 25.6005
R3835 VSS.n481 VSS.n269 25.6005
R3836 VSS.n487 VSS.n269 25.6005
R3837 VSS.n488 VSS.n487 25.6005
R3838 VSS.n489 VSS.n488 25.6005
R3839 VSS.n489 VSS.n267 25.6005
R3840 VSS.n495 VSS.n267 25.6005
R3841 VSS.n496 VSS.n495 25.6005
R3842 VSS.n497 VSS.n496 25.6005
R3843 VSS.n497 VSS.n265 25.6005
R3844 VSS.n503 VSS.n265 25.6005
R3845 VSS.n504 VSS.n503 25.6005
R3846 VSS.n505 VSS.n504 25.6005
R3847 VSS.n505 VSS.n263 25.6005
R3848 VSS.n511 VSS.n263 25.6005
R3849 VSS.n512 VSS.n511 25.6005
R3850 VSS.n513 VSS.n255 25.6005
R3851 VSS.n523 VSS.n255 25.6005
R3852 VSS.n524 VSS.n523 25.6005
R3853 VSS.n525 VSS.n524 25.6005
R3854 VSS.n525 VSS.n248 25.6005
R3855 VSS.n2298 VSS.n248 25.6005
R3856 VSS.n2299 VSS.n2298 25.6005
R3857 VSS.n2300 VSS.n2299 25.6005
R3858 VSS.n2300 VSS.n241 25.6005
R3859 VSS.n2311 VSS.n241 25.6005
R3860 VSS.n2312 VSS.n2311 25.6005
R3861 VSS.n2313 VSS.n2312 25.6005
R3862 VSS.n2313 VSS.n234 25.6005
R3863 VSS.n2324 VSS.n234 25.6005
R3864 VSS.n2325 VSS.n2324 25.6005
R3865 VSS.n2326 VSS.n2325 25.6005
R3866 VSS.n2326 VSS.n227 25.6005
R3867 VSS.n2337 VSS.n227 25.6005
R3868 VSS.n2338 VSS.n2337 25.6005
R3869 VSS.n2339 VSS.n2338 25.6005
R3870 VSS.n2339 VSS.n220 25.6005
R3871 VSS.n2350 VSS.n220 25.6005
R3872 VSS.n2351 VSS.n2350 25.6005
R3873 VSS.n2352 VSS.n2351 25.6005
R3874 VSS.n2352 VSS.n212 25.6005
R3875 VSS.n2362 VSS.n212 25.6005
R3876 VSS.n2363 VSS.n2362 25.6005
R3877 VSS.n2364 VSS.n2363 25.6005
R3878 VSS.n2364 VSS.n204 25.6005
R3879 VSS.n2374 VSS.n204 25.6005
R3880 VSS.n2375 VSS.n2374 25.6005
R3881 VSS.n2376 VSS.n2375 25.6005
R3882 VSS.n2376 VSS.n196 25.6005
R3883 VSS.n2386 VSS.n196 25.6005
R3884 VSS.n2387 VSS.n2386 25.6005
R3885 VSS.n2388 VSS.n2387 25.6005
R3886 VSS.n2388 VSS.n187 25.6005
R3887 VSS.n2398 VSS.n187 25.6005
R3888 VSS.n2399 VSS.n2398 25.6005
R3889 VSS.n2400 VSS.n2399 25.6005
R3890 VSS.n2400 VSS.n179 25.6005
R3891 VSS.n2410 VSS.n179 25.6005
R3892 VSS.n2411 VSS.n2410 25.6005
R3893 VSS.n2412 VSS.n2411 25.6005
R3894 VSS.n2412 VSS.n171 25.6005
R3895 VSS.n2422 VSS.n171 25.6005
R3896 VSS.n2423 VSS.n2422 25.6005
R3897 VSS.n2424 VSS.n2423 25.6005
R3898 VSS.n2424 VSS.n163 25.6005
R3899 VSS.n2434 VSS.n163 25.6005
R3900 VSS.n2435 VSS.n2434 25.6005
R3901 VSS.n2436 VSS.n2435 25.6005
R3902 VSS.n2436 VSS.n155 25.6005
R3903 VSS.n2446 VSS.n155 25.6005
R3904 VSS.n2447 VSS.n2446 25.6005
R3905 VSS.n2448 VSS.n2447 25.6005
R3906 VSS.n2448 VSS.n148 25.6005
R3907 VSS.n2458 VSS.n148 25.6005
R3908 VSS.n2459 VSS.n2458 25.6005
R3909 VSS.n2487 VSS.n2459 25.6005
R3910 VSS.n2487 VSS.n2486 25.6005
R3911 VSS.n2539 VSS.n2538 25.6005
R3912 VSS.n2538 VSS.n2537 25.6005
R3913 VSS.n2537 VSS.n2536 25.6005
R3914 VSS.n2536 VSS.n2534 25.6005
R3915 VSS.n2534 VSS.n2531 25.6005
R3916 VSS.n2531 VSS.n2530 25.6005
R3917 VSS.n2530 VSS.n2527 25.6005
R3918 VSS.n2527 VSS.n2526 25.6005
R3919 VSS.n2526 VSS.n2523 25.6005
R3920 VSS.n2523 VSS.n2522 25.6005
R3921 VSS.n2522 VSS.n2519 25.6005
R3922 VSS.n2519 VSS.n2518 25.6005
R3923 VSS.n2518 VSS.n2515 25.6005
R3924 VSS.n2515 VSS.n2514 25.6005
R3925 VSS.n2514 VSS.n2511 25.6005
R3926 VSS.n2511 VSS.n2510 25.6005
R3927 VSS.n2510 VSS.n2507 25.6005
R3928 VSS.n2507 VSS.n2506 25.6005
R3929 VSS.n2506 VSS.n2503 25.6005
R3930 VSS.n2496 VSS.n2493 25.6005
R3931 VSS.n2545 VSS.n117 25.6005
R3932 VSS.n2545 VSS.n118 25.6005
R3933 VSS.n2460 VSS.n118 25.6005
R3934 VSS.n2463 VSS.n2460 25.6005
R3935 VSS.n2464 VSS.n2463 25.6005
R3936 VSS.n2467 VSS.n2464 25.6005
R3937 VSS.n2468 VSS.n2467 25.6005
R3938 VSS.n2471 VSS.n2468 25.6005
R3939 VSS.n2472 VSS.n2471 25.6005
R3940 VSS.n2475 VSS.n2472 25.6005
R3941 VSS.n2476 VSS.n2475 25.6005
R3942 VSS.n2479 VSS.n2476 25.6005
R3943 VSS.n2480 VSS.n2479 25.6005
R3944 VSS.n2483 VSS.n2480 25.6005
R3945 VSS.n2485 VSS.n2483 25.6005
R3946 VSS.n1801 VSS.n855 25.6005
R3947 VSS.n1802 VSS.n1801 25.6005
R3948 VSS.n1803 VSS.n1802 25.6005
R3949 VSS.n1803 VSS.n829 25.6005
R3950 VSS.n1876 VSS.n829 25.6005
R3951 VSS.n1876 VSS.n1875 25.6005
R3952 VSS.n1875 VSS.n1874 25.6005
R3953 VSS.n1874 VSS.n1873 25.6005
R3954 VSS.n1873 VSS.n830 25.6005
R3955 VSS.n837 VSS.n830 25.6005
R3956 VSS.n1866 VSS.n837 25.6005
R3957 VSS.n1785 VSS.n1784 25.6005
R3958 VSS.n1784 VSS.n1783 25.6005
R3959 VSS.n1783 VSS.n1780 25.6005
R3960 VSS.n1780 VSS.n1779 25.6005
R3961 VSS.n1779 VSS.n1776 25.6005
R3962 VSS.n1776 VSS.n1775 25.6005
R3963 VSS.n1775 VSS.n1772 25.6005
R3964 VSS.n1772 VSS.n1771 25.6005
R3965 VSS.n1771 VSS.n1768 25.6005
R3966 VSS.n1768 VSS.n1767 25.6005
R3967 VSS.n1767 VSS.n1764 25.6005
R3968 VSS.n1764 VSS.n1763 25.6005
R3969 VSS.n1763 VSS.n1760 25.6005
R3970 VSS.n1760 VSS.n1759 25.6005
R3971 VSS.n1759 VSS.n1756 25.6005
R3972 VSS.n1756 VSS.n1755 25.6005
R3973 VSS.n1755 VSS.n1752 25.6005
R3974 VSS.n1752 VSS.n1751 25.6005
R3975 VSS.n1751 VSS.n1748 25.6005
R3976 VSS.n1748 VSS.n1747 25.6005
R3977 VSS.n1747 VSS.n1744 25.6005
R3978 VSS.n1744 VSS.n1743 25.6005
R3979 VSS.n1739 VSS.n1738 25.6005
R3980 VSS.n1738 VSS.n1737 25.6005
R3981 VSS.n1737 VSS.n850 25.6005
R3982 VSS.n1809 VSS.n850 25.6005
R3983 VSS.n1810 VSS.n1809 25.6005
R3984 VSS.n1812 VSS.n1810 25.6005
R3985 VSS.n1813 VSS.n1812 25.6005
R3986 VSS.n1815 VSS.n1813 25.6005
R3987 VSS.n1816 VSS.n1815 25.6005
R3988 VSS.n1817 VSS.n1816 25.6005
R3989 VSS.n1818 VSS.n1817 25.6005
R3990 VSS.n1865 VSS.n1864 25.6005
R3991 VSS.n1864 VSS.n838 25.6005
R3992 VSS.n1859 VSS.n838 25.6005
R3993 VSS.n1859 VSS.n1858 25.6005
R3994 VSS.n1858 VSS.n840 25.6005
R3995 VSS.n1853 VSS.n840 25.6005
R3996 VSS.n1853 VSS.n1852 25.6005
R3997 VSS.n1852 VSS.n1851 25.6005
R3998 VSS.n1851 VSS.n842 25.6005
R3999 VSS.n1842 VSS.n1841 25.6005
R4000 VSS.n1841 VSS.n845 25.6005
R4001 VSS.n1835 VSS.n845 25.6005
R4002 VSS.n1835 VSS.n1834 25.6005
R4003 VSS.n1834 VSS.n1833 25.6005
R4004 VSS.n1833 VSS.n847 25.6005
R4005 VSS.n1827 VSS.n847 25.6005
R4006 VSS.n1827 VSS.n1826 25.6005
R4007 VSS.n1826 VSS.n1825 25.6005
R4008 VSS.n1825 VSS.n849 25.6005
R4009 VSS.n1819 VSS.n849 25.6005
R4010 VSS.n1292 VSS.n1229 25.6005
R4011 VSS.n1326 VSS.n1229 25.6005
R4012 VSS.n1326 VSS.n1325 25.6005
R4013 VSS.n1325 VSS.n1324 25.6005
R4014 VSS.n1324 VSS.n1230 25.6005
R4015 VSS.n1307 VSS.n1230 25.6005
R4016 VSS.n1307 VSS.n1104 25.6005
R4017 VSS.n1532 VSS.n1104 25.6005
R4018 VSS.n1533 VSS.n1532 25.6005
R4019 VSS.n1534 VSS.n1533 25.6005
R4020 VSS.n1534 VSS.n1094 25.6005
R4021 VSS.n1291 VSS.n1290 25.6005
R4022 VSS.n1290 VSS.n1237 25.6005
R4023 VSS.n1238 VSS.n1237 25.6005
R4024 VSS.n1283 VSS.n1238 25.6005
R4025 VSS.n1283 VSS.n1282 25.6005
R4026 VSS.n1282 VSS.n1281 25.6005
R4027 VSS.n1281 VSS.n1240 25.6005
R4028 VSS.n1276 VSS.n1240 25.6005
R4029 VSS.n1276 VSS.n1275 25.6005
R4030 VSS.n1275 VSS.n1274 25.6005
R4031 VSS.n1274 VSS.n1243 25.6005
R4032 VSS.n1269 VSS.n1243 25.6005
R4033 VSS.n1269 VSS.n1268 25.6005
R4034 VSS.n1268 VSS.n1267 25.6005
R4035 VSS.n1267 VSS.n1246 25.6005
R4036 VSS.n1262 VSS.n1246 25.6005
R4037 VSS.n1262 VSS.n1261 25.6005
R4038 VSS.n1261 VSS.n1260 25.6005
R4039 VSS.n1260 VSS.n1249 25.6005
R4040 VSS.n1255 VSS.n1249 25.6005
R4041 VSS.n1255 VSS.n1254 25.6005
R4042 VSS.n1254 VSS.n1253 25.6005
R4043 VSS.n1297 VSS.n1234 25.6005
R4044 VSS.n1298 VSS.n1297 25.6005
R4045 VSS.n1301 VSS.n1298 25.6005
R4046 VSS.n1302 VSS.n1301 25.6005
R4047 VSS.n1303 VSS.n1302 25.6005
R4048 VSS.n1303 VSS.n1108 25.6005
R4049 VSS.n1521 VSS.n1108 25.6005
R4050 VSS.n1522 VSS.n1521 25.6005
R4051 VSS.n1526 VSS.n1525 25.6005
R4052 VSS.n1588 VSS.n1587 25.6005
R4053 VSS.n1587 VSS.n1586 25.6005
R4054 VSS.n1586 VSS.n1585 25.6005
R4055 VSS.n1585 VSS.n1583 25.6005
R4056 VSS.n1583 VSS.n1580 25.6005
R4057 VSS.n1580 VSS.n1579 25.6005
R4058 VSS.n1579 VSS.n1576 25.6005
R4059 VSS.n1576 VSS.n1575 25.6005
R4060 VSS.n1575 VSS.n1572 25.6005
R4061 VSS.n1572 VSS.n1571 25.6005
R4062 VSS.n1571 VSS.n1568 25.6005
R4063 VSS.n1568 VSS.n1567 25.6005
R4064 VSS.n1567 VSS.n1564 25.6005
R4065 VSS.n1564 VSS.n1563 25.6005
R4066 VSS.n1563 VSS.n1560 25.6005
R4067 VSS.n1560 VSS.n1559 25.6005
R4068 VSS.n1559 VSS.n1556 25.6005
R4069 VSS.n1556 VSS.n1555 25.6005
R4070 VSS.n1555 VSS.n1552 25.6005
R4071 VSS.n1552 VSS.n1551 25.6005
R4072 VSS.n1551 VSS.n1548 25.6005
R4073 VSS.n1548 VSS.n1547 25.6005
R4074 VSS.n1468 VSS.n1467 25.6005
R4075 VSS.n1469 VSS.n1468 25.6005
R4076 VSS.n1469 VSS.n1115 25.6005
R4077 VSS.n1475 VSS.n1115 25.6005
R4078 VSS.n1476 VSS.n1475 25.6005
R4079 VSS.n1516 VSS.n1476 25.6005
R4080 VSS.n1516 VSS.n1515 25.6005
R4081 VSS.n1515 VSS.n1514 25.6005
R4082 VSS.n1514 VSS.n1477 25.6005
R4083 VSS.n1509 VSS.n1477 25.6005
R4084 VSS.n1509 VSS.n1508 25.6005
R4085 VSS.n1508 VSS.n1507 25.6005
R4086 VSS.n1507 VSS.n1479 25.6005
R4087 VSS.n1481 VSS.n1479 25.6005
R4088 VSS.n1483 VSS.n1481 25.6005
R4089 VSS.n1496 VSS.n1495 25.6005
R4090 VSS.n1492 VSS.n1485 25.6005
R4091 VSS.n1486 VSS.n1485 25.6005
R4092 VSS.n1486 VSS.n749 25.6005
R4093 VSS.n2094 VSS.n754 25.6005
R4094 VSS.n2094 VSS.n2093 25.6005
R4095 VSS.n2093 VSS.n2092 25.6005
R4096 VSS.n2092 VSS.n755 25.6005
R4097 VSS.n2086 VSS.n755 25.6005
R4098 VSS.n2086 VSS.n2085 25.6005
R4099 VSS.n2085 VSS.n2084 25.6005
R4100 VSS.n2084 VSS.n759 25.6005
R4101 VSS.n2078 VSS.n759 25.6005
R4102 VSS.n2078 VSS.n2077 25.6005
R4103 VSS.n2077 VSS.n2076 25.6005
R4104 VSS.n2076 VSS.n763 25.6005
R4105 VSS.n2070 VSS.n763 25.6005
R4106 VSS.n2070 VSS.n2069 25.6005
R4107 VSS.n2069 VSS.n2068 25.6005
R4108 VSS.n1131 VSS.n1118 25.6005
R4109 VSS.n1134 VSS.n1131 25.6005
R4110 VSS.n1135 VSS.n1134 25.6005
R4111 VSS.n1138 VSS.n1135 25.6005
R4112 VSS.n1139 VSS.n1138 25.6005
R4113 VSS.n1142 VSS.n1139 25.6005
R4114 VSS.n1143 VSS.n1142 25.6005
R4115 VSS.n1146 VSS.n1143 25.6005
R4116 VSS.n1147 VSS.n1146 25.6005
R4117 VSS.n1150 VSS.n1147 25.6005
R4118 VSS.n1151 VSS.n1150 25.6005
R4119 VSS.n1154 VSS.n1151 25.6005
R4120 VSS.n1155 VSS.n1154 25.6005
R4121 VSS.n1158 VSS.n1155 25.6005
R4122 VSS.n1159 VSS.n1158 25.6005
R4123 VSS.n1162 VSS.n1159 25.6005
R4124 VSS.n1164 VSS.n1162 25.6005
R4125 VSS.n1165 VSS.n1164 25.6005
R4126 VSS.n1460 VSS.n1165 25.6005
R4127 VSS.n1460 VSS.n1459 25.6005
R4128 VSS.n1459 VSS.n1458 25.6005
R4129 VSS.n1458 VSS.n1166 25.6005
R4130 VSS.n1453 VSS.n1452 25.6005
R4131 VSS.n1452 VSS.n1451 25.6005
R4132 VSS.n1451 VSS.n1170 25.6005
R4133 VSS.n1446 VSS.n1170 25.6005
R4134 VSS.n1446 VSS.n1445 25.6005
R4135 VSS.n1445 VSS.n1444 25.6005
R4136 VSS.n1444 VSS.n1173 25.6005
R4137 VSS.n1439 VSS.n1173 25.6005
R4138 VSS.n1439 VSS.n1438 25.6005
R4139 VSS.n1438 VSS.n1437 25.6005
R4140 VSS.n1437 VSS.n1176 25.6005
R4141 VSS.n1432 VSS.n1176 25.6005
R4142 VSS.n1432 VSS.n1431 25.6005
R4143 VSS.n1431 VSS.n1430 25.6005
R4144 VSS.n1430 VSS.n1179 25.6005
R4145 VSS.n1425 VSS.n1179 25.6005
R4146 VSS.n1425 VSS.n1424 25.6005
R4147 VSS.n1424 VSS.n1423 25.6005
R4148 VSS.n1423 VSS.n1182 25.6005
R4149 VSS.n1418 VSS.n1182 25.6005
R4150 VSS.n1418 VSS.n1417 25.6005
R4151 VSS.n1417 VSS.n1416 25.6005
R4152 VSS.n1416 VSS.n1185 25.6005
R4153 VSS.n1411 VSS.n1410 25.6005
R4154 VSS.n1410 VSS.n1409 25.6005
R4155 VSS.n1409 VSS.n1188 25.6005
R4156 VSS.n1404 VSS.n1188 25.6005
R4157 VSS.n1404 VSS.n1403 25.6005
R4158 VSS.n1403 VSS.n1402 25.6005
R4159 VSS.n1402 VSS.n1191 25.6005
R4160 VSS.n1397 VSS.n1191 25.6005
R4161 VSS.n1397 VSS.n1396 25.6005
R4162 VSS.n1396 VSS.n1395 25.6005
R4163 VSS.n1395 VSS.n1194 25.6005
R4164 VSS.n1390 VSS.n1194 25.6005
R4165 VSS.n1390 VSS.n1389 25.6005
R4166 VSS.n1389 VSS.n1388 25.6005
R4167 VSS.n1388 VSS.n1197 25.6005
R4168 VSS.n1383 VSS.n1197 25.6005
R4169 VSS.n1383 VSS.n1382 25.6005
R4170 VSS.n1382 VSS.n1381 25.6005
R4171 VSS.n1381 VSS.n1200 25.6005
R4172 VSS.n1376 VSS.n1200 25.6005
R4173 VSS.n1376 VSS.n1375 25.6005
R4174 VSS.n1375 VSS.n1374 25.6005
R4175 VSS.n1374 VSS.n1203 25.6005
R4176 VSS.n1369 VSS.n1368 25.6005
R4177 VSS.n1368 VSS.n1367 25.6005
R4178 VSS.n1367 VSS.n1206 25.6005
R4179 VSS.n1362 VSS.n1206 25.6005
R4180 VSS.n1362 VSS.n1361 25.6005
R4181 VSS.n1361 VSS.n1360 25.6005
R4182 VSS.n1360 VSS.n1209 25.6005
R4183 VSS.n1355 VSS.n1209 25.6005
R4184 VSS.n1355 VSS.n1354 25.6005
R4185 VSS.n1354 VSS.n1353 25.6005
R4186 VSS.n1353 VSS.n1212 25.6005
R4187 VSS.n1348 VSS.n1212 25.6005
R4188 VSS.n1348 VSS.n1347 25.6005
R4189 VSS.n1347 VSS.n1346 25.6005
R4190 VSS.n1346 VSS.n1215 25.6005
R4191 VSS.n1341 VSS.n1215 25.6005
R4192 VSS.n1341 VSS.n1340 25.6005
R4193 VSS.n1340 VSS.n1339 25.6005
R4194 VSS.n1339 VSS.n1218 25.6005
R4195 VSS.n1334 VSS.n1218 25.6005
R4196 VSS.n1334 VSS.n1333 25.6005
R4197 VSS.n1333 VSS.n1332 25.6005
R4198 VSS.n1312 VSS.n1221 25.6005
R4199 VSS.n1313 VSS.n1312 25.6005
R4200 VSS.n1319 VSS.n1313 25.6005
R4201 VSS.n1319 VSS.n1318 25.6005
R4202 VSS.n1318 VSS.n1317 25.6005
R4203 VSS.n1317 VSS.n1314 25.6005
R4204 VSS.n1314 VSS.n1101 25.6005
R4205 VSS.n1539 VSS.n1101 25.6005
R4206 VSS.n1540 VSS.n1539 25.6005
R4207 VSS.n1541 VSS.n1540 25.6005
R4208 VSS.n1541 VSS.n1078 25.6005
R4209 VSS.n1595 VSS.n1078 25.6005
R4210 VSS.n1596 VSS.n1595 25.6005
R4211 VSS.n1598 VSS.n1596 25.6005
R4212 VSS.n1598 VSS.n1597 25.6005
R4213 VSS.n1619 VSS.n1013 25.6005
R4214 VSS.n1634 VSS.n910 25.6005
R4215 VSS.n1634 VSS.n1633 25.6005
R4216 VSS.n1633 VSS.n1632 25.6005
R4217 VSS.n1665 VSS.n888 25.6005
R4218 VSS.n1666 VSS.n1665 25.6005
R4219 VSS.n1667 VSS.n1666 25.6005
R4220 VSS.n1667 VSS.n866 25.6005
R4221 VSS.n1720 VSS.n866 25.6005
R4222 VSS.n1721 VSS.n1720 25.6005
R4223 VSS.n1722 VSS.n1721 25.6005
R4224 VSS.n1722 VSS.n862 25.6005
R4225 VSS.n1791 VSS.n862 25.6005
R4226 VSS.n1792 VSS.n1791 25.6005
R4227 VSS.n1796 VSS.n1792 25.6005
R4228 VSS.n1796 VSS.n1795 25.6005
R4229 VSS.n1795 VSS.n1794 25.6005
R4230 VSS.n1794 VSS.n823 25.6005
R4231 VSS.n1881 VSS.n823 25.6005
R4232 VSS.n2062 VSS.n767 25.6005
R4233 VSS.n2062 VSS.n2061 25.6005
R4234 VSS.n2061 VSS.n2060 25.6005
R4235 VSS.n2060 VSS.n2058 25.6005
R4236 VSS.n2058 VSS.n2055 25.6005
R4237 VSS.n2055 VSS.n2054 25.6005
R4238 VSS.n2054 VSS.n2051 25.6005
R4239 VSS.n2051 VSS.n2050 25.6005
R4240 VSS.n2050 VSS.n2047 25.6005
R4241 VSS.n2047 VSS.n2046 25.6005
R4242 VSS.n2046 VSS.n2043 25.6005
R4243 VSS.n2043 VSS.n2042 25.6005
R4244 VSS.n2042 VSS.n2039 25.6005
R4245 VSS.n2039 VSS.n2038 25.6005
R4246 VSS.n2038 VSS.n2035 25.6005
R4247 VSS.n2035 VSS.n2034 25.6005
R4248 VSS.n2034 VSS.n2031 25.6005
R4249 VSS.n2031 VSS.n2030 25.6005
R4250 VSS.n2030 VSS.n2028 25.6005
R4251 VSS.n2028 VSS.n2027 25.6005
R4252 VSS.n2027 VSS.n780 25.6005
R4253 VSS.n2022 VSS.n780 25.6005
R4254 VSS.n2021 VSS.n2020 25.6005
R4255 VSS.n2020 VSS.n2017 25.6005
R4256 VSS.n2017 VSS.n2016 25.6005
R4257 VSS.n2016 VSS.n2013 25.6005
R4258 VSS.n2013 VSS.n2012 25.6005
R4259 VSS.n2012 VSS.n2009 25.6005
R4260 VSS.n2009 VSS.n2008 25.6005
R4261 VSS.n2008 VSS.n2005 25.6005
R4262 VSS.n2005 VSS.n2004 25.6005
R4263 VSS.n2004 VSS.n2001 25.6005
R4264 VSS.n2001 VSS.n2000 25.6005
R4265 VSS.n2000 VSS.n1997 25.6005
R4266 VSS.n1997 VSS.n1996 25.6005
R4267 VSS.n1996 VSS.n1993 25.6005
R4268 VSS.n1993 VSS.n1992 25.6005
R4269 VSS.n1992 VSS.n1989 25.6005
R4270 VSS.n1989 VSS.n1988 25.6005
R4271 VSS.n1988 VSS.n1985 25.6005
R4272 VSS.n1985 VSS.n1984 25.6005
R4273 VSS.n1984 VSS.n1981 25.6005
R4274 VSS.n1981 VSS.n1980 25.6005
R4275 VSS.n1980 VSS.n1977 25.6005
R4276 VSS.n1977 VSS.n1976 25.6005
R4277 VSS.n1973 VSS.n1972 25.6005
R4278 VSS.n1972 VSS.n1969 25.6005
R4279 VSS.n1969 VSS.n1968 25.6005
R4280 VSS.n1968 VSS.n1965 25.6005
R4281 VSS.n1965 VSS.n1964 25.6005
R4282 VSS.n1964 VSS.n1961 25.6005
R4283 VSS.n1961 VSS.n1960 25.6005
R4284 VSS.n1960 VSS.n1957 25.6005
R4285 VSS.n1957 VSS.n1956 25.6005
R4286 VSS.n1956 VSS.n1953 25.6005
R4287 VSS.n1953 VSS.n1952 25.6005
R4288 VSS.n1952 VSS.n1949 25.6005
R4289 VSS.n1949 VSS.n1948 25.6005
R4290 VSS.n1948 VSS.n1945 25.6005
R4291 VSS.n1945 VSS.n1944 25.6005
R4292 VSS.n1944 VSS.n1941 25.6005
R4293 VSS.n1941 VSS.n1940 25.6005
R4294 VSS.n1940 VSS.n1937 25.6005
R4295 VSS.n1937 VSS.n1936 25.6005
R4296 VSS.n1936 VSS.n1933 25.6005
R4297 VSS.n1933 VSS.n1932 25.6005
R4298 VSS.n1932 VSS.n1929 25.6005
R4299 VSS.n1929 VSS.n1928 25.6005
R4300 VSS.n1925 VSS.n1924 25.6005
R4301 VSS.n1924 VSS.n1921 25.6005
R4302 VSS.n1921 VSS.n1920 25.6005
R4303 VSS.n1920 VSS.n1917 25.6005
R4304 VSS.n1917 VSS.n1916 25.6005
R4305 VSS.n1916 VSS.n1913 25.6005
R4306 VSS.n1913 VSS.n1912 25.6005
R4307 VSS.n1912 VSS.n1909 25.6005
R4308 VSS.n1909 VSS.n1908 25.6005
R4309 VSS.n1908 VSS.n1905 25.6005
R4310 VSS.n1905 VSS.n1904 25.6005
R4311 VSS.n1904 VSS.n1901 25.6005
R4312 VSS.n1901 VSS.n1900 25.6005
R4313 VSS.n1900 VSS.n1897 25.6005
R4314 VSS.n1897 VSS.n1896 25.6005
R4315 VSS.n1896 VSS.n1893 25.6005
R4316 VSS.n1893 VSS.n1892 25.6005
R4317 VSS.n1892 VSS.n1889 25.6005
R4318 VSS.n1889 VSS.n1888 25.6005
R4319 VSS.n1888 VSS.n1885 25.6005
R4320 VSS.n1885 VSS.n1884 25.6005
R4321 VSS.n1884 VSS.n1882 25.6005
R4322 VSS.n2115 VSS.n2114 25.6005
R4323 VSS.n2114 VSS.n643 25.6005
R4324 VSS.n2109 VSS.n643 25.6005
R4325 VSS.n2116 VSS.n635 25.6005
R4326 VSS.n2126 VSS.n635 25.6005
R4327 VSS.n2127 VSS.n2126 25.6005
R4328 VSS.n2128 VSS.n2127 25.6005
R4329 VSS.n2128 VSS.n627 25.6005
R4330 VSS.n2138 VSS.n627 25.6005
R4331 VSS.n2139 VSS.n2138 25.6005
R4332 VSS.n2140 VSS.n2139 25.6005
R4333 VSS.n2140 VSS.n619 25.6005
R4334 VSS.n2150 VSS.n619 25.6005
R4335 VSS.n2151 VSS.n2150 25.6005
R4336 VSS.n2152 VSS.n2151 25.6005
R4337 VSS.n2152 VSS.n610 25.6005
R4338 VSS.n2162 VSS.n610 25.6005
R4339 VSS.n2163 VSS.n2162 25.6005
R4340 VSS.n2164 VSS.n2163 25.6005
R4341 VSS.n2164 VSS.n602 25.6005
R4342 VSS.n2174 VSS.n602 25.6005
R4343 VSS.n2175 VSS.n2174 25.6005
R4344 VSS.n2176 VSS.n2175 25.6005
R4345 VSS.n2176 VSS.n594 25.6005
R4346 VSS.n2186 VSS.n594 25.6005
R4347 VSS.n2187 VSS.n2186 25.6005
R4348 VSS.n2188 VSS.n2187 25.6005
R4349 VSS.n2188 VSS.n586 25.6005
R4350 VSS.n2198 VSS.n586 25.6005
R4351 VSS.n2199 VSS.n2198 25.6005
R4352 VSS.n2200 VSS.n2199 25.6005
R4353 VSS.n2200 VSS.n578 25.6005
R4354 VSS.n2210 VSS.n578 25.6005
R4355 VSS.n2211 VSS.n2210 25.6005
R4356 VSS.n2212 VSS.n2211 25.6005
R4357 VSS.n2212 VSS.n570 25.6005
R4358 VSS.n2222 VSS.n570 25.6005
R4359 VSS.n2223 VSS.n2222 25.6005
R4360 VSS.n2224 VSS.n2223 25.6005
R4361 VSS.n2224 VSS.n562 25.6005
R4362 VSS.n2234 VSS.n562 25.6005
R4363 VSS.n2235 VSS.n2234 25.6005
R4364 VSS.n2236 VSS.n2235 25.6005
R4365 VSS.n2236 VSS.n554 25.6005
R4366 VSS.n2246 VSS.n554 25.6005
R4367 VSS.n2247 VSS.n2246 25.6005
R4368 VSS.n2248 VSS.n2247 25.6005
R4369 VSS.n2248 VSS.n546 25.6005
R4370 VSS.n2258 VSS.n546 25.6005
R4371 VSS.n2259 VSS.n2258 25.6005
R4372 VSS.n2260 VSS.n2259 25.6005
R4373 VSS.n2260 VSS.n538 25.6005
R4374 VSS.n2271 VSS.n538 25.6005
R4375 VSS.n2272 VSS.n2271 25.6005
R4376 VSS.n2273 VSS.n2272 25.6005
R4377 VSS.n2273 VSS.n532 25.6005
R4378 VSS.n2285 VSS.n2284 25.6005
R4379 VSS.n2284 VSS.n2283 25.6005
R4380 VSS.n2283 VSS.n2280 25.6005
R4381 VSS.n2280 VSS.n2279 25.6005
R4382 VSS.n2121 VSS.n2120 25.6005
R4383 VSS.n2122 VSS.n2121 25.6005
R4384 VSS.n2122 VSS.n631 25.6005
R4385 VSS.n2132 VSS.n631 25.6005
R4386 VSS.n2133 VSS.n2132 25.6005
R4387 VSS.n2134 VSS.n2133 25.6005
R4388 VSS.n2134 VSS.n623 25.6005
R4389 VSS.n2144 VSS.n623 25.6005
R4390 VSS.n2145 VSS.n2144 25.6005
R4391 VSS.n2146 VSS.n2145 25.6005
R4392 VSS.n2146 VSS.n614 25.6005
R4393 VSS.n2156 VSS.n614 25.6005
R4394 VSS.n2157 VSS.n2156 25.6005
R4395 VSS.n2158 VSS.n2157 25.6005
R4396 VSS.n2158 VSS.n606 25.6005
R4397 VSS.n2168 VSS.n606 25.6005
R4398 VSS.n2169 VSS.n2168 25.6005
R4399 VSS.n2170 VSS.n2169 25.6005
R4400 VSS.n2170 VSS.n598 25.6005
R4401 VSS.n2180 VSS.n598 25.6005
R4402 VSS.n2181 VSS.n2180 25.6005
R4403 VSS.n2182 VSS.n2181 25.6005
R4404 VSS.n2182 VSS.n590 25.6005
R4405 VSS.n2192 VSS.n590 25.6005
R4406 VSS.n2193 VSS.n2192 25.6005
R4407 VSS.n2194 VSS.n2193 25.6005
R4408 VSS.n2194 VSS.n582 25.6005
R4409 VSS.n2204 VSS.n582 25.6005
R4410 VSS.n2205 VSS.n2204 25.6005
R4411 VSS.n2206 VSS.n2205 25.6005
R4412 VSS.n2206 VSS.n574 25.6005
R4413 VSS.n2216 VSS.n574 25.6005
R4414 VSS.n2217 VSS.n2216 25.6005
R4415 VSS.n2218 VSS.n2217 25.6005
R4416 VSS.n2218 VSS.n566 25.6005
R4417 VSS.n2228 VSS.n566 25.6005
R4418 VSS.n2229 VSS.n2228 25.6005
R4419 VSS.n2230 VSS.n2229 25.6005
R4420 VSS.n2230 VSS.n558 25.6005
R4421 VSS.n2240 VSS.n558 25.6005
R4422 VSS.n2241 VSS.n2240 25.6005
R4423 VSS.n2242 VSS.n2241 25.6005
R4424 VSS.n2242 VSS.n550 25.6005
R4425 VSS.n2252 VSS.n550 25.6005
R4426 VSS.n2253 VSS.n2252 25.6005
R4427 VSS.n2254 VSS.n2253 25.6005
R4428 VSS.n2254 VSS.n542 25.6005
R4429 VSS.n2264 VSS.n542 25.6005
R4430 VSS.n2265 VSS.n2264 25.6005
R4431 VSS.n2267 VSS.n2265 25.6005
R4432 VSS.n2267 VSS.n2266 25.6005
R4433 VSS.n2266 VSS.n535 25.6005
R4434 VSS.n535 VSS.n533 25.6005
R4435 VSS.n1605 VSS.n1604 25.6005
R4436 VSS.n1604 VSS.n1026 25.6005
R4437 VSS.n1038 VSS.n1026 25.6005
R4438 VSS.n1041 VSS.n1038 25.6005
R4439 VSS.n1042 VSS.n1041 25.6005
R4440 VSS.n1045 VSS.n1042 25.6005
R4441 VSS.n1046 VSS.n1045 25.6005
R4442 VSS.n1049 VSS.n1046 25.6005
R4443 VSS.n1050 VSS.n1049 25.6005
R4444 VSS.n1053 VSS.n1050 25.6005
R4445 VSS.n1054 VSS.n1053 25.6005
R4446 VSS.n1057 VSS.n1054 25.6005
R4447 VSS.n1058 VSS.n1057 25.6005
R4448 VSS.n1061 VSS.n1058 25.6005
R4449 VSS.n1062 VSS.n1061 25.6005
R4450 VSS.n1065 VSS.n1062 25.6005
R4451 VSS.n1066 VSS.n1065 25.6005
R4452 VSS.n1069 VSS.n1066 25.6005
R4453 VSS.n1071 VSS.n1069 25.6005
R4454 VSS.n1072 VSS.n1071 25.6005
R4455 VSS.n1073 VSS.n1072 25.6005
R4456 VSS.n1073 VSS.n1019 25.6005
R4457 VSS.n1607 VSS.n1606 25.6005
R4458 VSS.n1606 VSS.n903 25.6005
R4459 VSS.n1639 VSS.n903 25.6005
R4460 VSS.n1640 VSS.n1639 25.6005
R4461 VSS.n1641 VSS.n1640 25.6005
R4462 VSS.n1641 VSS.n894 25.6005
R4463 VSS.n1657 VSS.n894 25.6005
R4464 VSS.n1658 VSS.n1657 25.6005
R4465 VSS.n1660 VSS.n1658 25.6005
R4466 VSS.n1660 VSS.n1659 25.6005
R4467 VSS.n1659 VSS.n882 25.6005
R4468 VSS.n1714 VSS.n1713 25.6005
R4469 VSS.n1713 VSS.n1712 25.6005
R4470 VSS.n1712 VSS.n1711 25.6005
R4471 VSS.n1711 VSS.n1709 25.6005
R4472 VSS.n1709 VSS.n1706 25.6005
R4473 VSS.n1706 VSS.n1705 25.6005
R4474 VSS.n1705 VSS.n1702 25.6005
R4475 VSS.n1702 VSS.n1701 25.6005
R4476 VSS.n1701 VSS.n1698 25.6005
R4477 VSS.n1698 VSS.n1697 25.6005
R4478 VSS.n1697 VSS.n1694 25.6005
R4479 VSS.n1694 VSS.n1693 25.6005
R4480 VSS.n1693 VSS.n1690 25.6005
R4481 VSS.n1690 VSS.n1689 25.6005
R4482 VSS.n1689 VSS.n1686 25.6005
R4483 VSS.n1686 VSS.n1685 25.6005
R4484 VSS.n1685 VSS.n1682 25.6005
R4485 VSS.n1682 VSS.n1681 25.6005
R4486 VSS.n1681 VSS.n1678 25.6005
R4487 VSS.n1678 VSS.n1677 25.6005
R4488 VSS.n1677 VSS.n1674 25.6005
R4489 VSS.n1674 VSS.n1673 25.6005
R4490 VSS.n1612 VSS.n1611 25.6005
R4491 VSS.n1614 VSS.n1612 25.6005
R4492 VSS.n1614 VSS.n1613 25.6005
R4493 VSS.n1613 VSS.n899 25.6005
R4494 VSS.n1645 VSS.n899 25.6005
R4495 VSS.n1646 VSS.n1645 25.6005
R4496 VSS.n1652 VSS.n1646 25.6005
R4497 VSS.n1648 VSS.n1647 25.6005
R4498 VSS.n1647 VSS.n883 25.6005
R4499 VSS.t91 VSS.n1869 25.0064
R4500 VSS.n351 VSS.n345 24.8476
R4501 VSS.n449 VSS.n443 24.8476
R4502 VSS.n421 VSS.n334 24.8476
R4503 VSS.n419 VSS.n332 24.8476
R4504 VSS.n5 VSS.n4 24.8476
R4505 VSS.n106 VSS.n88 24.8476
R4506 VSS.n60 VSS.n59 24.8476
R4507 VSS.n326 VSS.n271 24.8476
R4508 VSS.n2500 VSS.n2499 24.8476
R4509 VSS.n1524 VSS.n1095 24.8476
R4510 VSS.n994 VSS.n964 24.8476
R4511 VSS.n933 VSS.n930 24.8476
R4512 VSS.n732 VSS.n731 24.8476
R4513 VSS.n671 VSS.n667 24.8476
R4514 VSS.n2101 VSS.n2100 24.8476
R4515 VSS.n1627 VSS.n1011 24.8476
R4516 VSS.n101 VSS.n100 24.75
R4517 VSS.n64 VSS.n63 24.75
R4518 VSS.n364 VSS.n340 24.2609
R4519 VSS.n358 VSS.n338 24.2609
R4520 VSS.n462 VSS.n456 24.2609
R4521 VSS.n467 VSS.n458 24.2609
R4522 VSS.n94 VSS.n90 24.2609
R4523 VSS.n68 VSS.n47 24.2609
R4524 VSS.n645 VSS.n639 23.7181
R4525 VSS.n1593 VSS.n1591 23.4436
R4526 VSS.n364 VSS.n341 23.3417
R4527 VSS.n358 VSS.n339 23.3417
R4528 VSS.n348 VSS.n344 23.3417
R4529 VSS.n462 VSS.n457 23.3417
R4530 VSS.n467 VSS.n459 23.3417
R4531 VSS.n446 VSS.n442 23.3417
R4532 VSS.n423 VSS.n335 23.3417
R4533 VSS.n417 VSS.n331 23.3417
R4534 VSS.n14 VSS.n6 23.3417
R4535 VSS.n110 VSS.n109 23.3417
R4536 VSS.n94 VSS.n91 23.3417
R4537 VSS.n69 VSS.n68 23.3417
R4538 VSS.n56 VSS.n51 23.3417
R4539 VSS.n993 VSS.n966 23.3417
R4540 VSS.n937 VSS.n936 23.3417
R4541 VSS.n728 VSS.n702 23.3417
R4542 VSS.n672 VSS.n665 23.3417
R4543 VSS.n1799 VSS.n857 22.9226
R4544 VSS.n1805 VSS.n852 22.9226
R4545 VSS.n1878 VSS.n825 22.9226
R4546 VSS.n1484 VSS.n1483 22.5887
R4547 VSS.n1597 VSS.n1012 22.5887
R4548 VSS.n1504 VSS.t0 22.5151
R4549 VSS.n757 VSS.t45 22.5151
R4550 VSS.n352 VSS.n351 22.4252
R4551 VSS.n450 VSS.n449 22.4252
R4552 VSS.n2302 VSS.t16 22.4016
R4553 VSS.n2438 VSS.t13 22.4016
R4554 VSS.n1494 VSS.n1492 22.2123
R4555 VSS.n1620 VSS.n910 22.2123
R4556 VSS.n31 VSS.n30 22.0256
R4557 VSS.n368 VSS.n367 21.8358
R4558 VSS.n371 VSS.n337 21.8358
R4559 VSS.n354 VSS.n343 21.8358
R4560 VSS.n474 VSS.n455 21.8358
R4561 VSS.n471 VSS.n470 21.8358
R4562 VSS.n452 VSS.n441 21.8358
R4563 VSS.n427 VSS.n426 21.8358
R4564 VSS.n415 VSS.n330 21.8358
R4565 VSS.n16 VSS.n7 21.8358
R4566 VSS.n112 VSS.n86 21.8358
R4567 VSS.n98 VSS.n97 21.8358
R4568 VSS.n71 VSS.n46 21.8358
R4569 VSS.n55 VSS.n52 21.8358
R4570 VSS.n1523 VSS.n1522 21.8358
R4571 VSS.n990 VSS.n989 21.8358
R4572 VSS.n940 VSS.n928 21.8358
R4573 VSS.n727 VSS.n704 21.8358
R4574 VSS.n676 VSS.n675 21.8358
R4575 VSS.n2366 VSS.t42 21.3597
R4576 VSS.t26 VSS.n198 21.3597
R4577 VSS.n480 VSS.n271 21.0829
R4578 VSS.n2499 VSS.n2497 21.0829
R4579 VSS.t1 VSS.n1518 20.3709
R4580 VSS.n2080 VSS.t5 20.3709
R4581 VSS.n18 VSS.n8 20.3299
R4582 VSS.n986 VSS.n968 20.3299
R4583 VSS.n941 VSS.n926 20.3299
R4584 VSS.n724 VSS.n723 20.3299
R4585 VSS.n679 VSS.n663 20.3299
R4586 VSS.n2322 VSS.t54 20.3178
R4587 VSS.n174 VSS.t84 20.3178
R4588 VSS.n1807 VSS.t8 20.3178
R4589 VSS.n319 VSS.n272 19.9534
R4590 VSS.n2503 VSS.n2502 19.9534
R4591 VSS.n1609 VSS.n1021 19.7969
R4592 VSS.n1024 VSS.n1022 19.7969
R4593 VSS.n1637 VSS.n905 19.7969
R4594 VSS.n1636 VSS.n907 19.7969
R4595 VSS.n1643 VSS.n901 19.7969
R4596 VSS.n1655 VSS.n896 19.7969
R4597 VSS.n1654 VSS.n890 19.7969
R4598 VSS.n1663 VSS.n1662 19.7969
R4599 VSS.n886 VSS.n885 19.7969
R4600 VSS.n1670 VSS.n1669 19.7969
R4601 VSS.n20 VSS.n9 18.824
R4602 VSS.n985 VSS.n970 18.824
R4603 VSS.n945 VSS.n944 18.824
R4604 VSS.n720 VSS.n706 18.824
R4605 VSS.n680 VSS.n661 18.824
R4606 VSS.n1329 VSS.n1224 18.7549
R4607 VSS.n1328 VSS.n1226 18.7549
R4608 VSS.n1322 VSS.n1321 18.7549
R4609 VSS.n1309 VSS.n1110 18.7549
R4610 VSS.n1530 VSS.n1529 18.7549
R4611 VSS.n1536 VSS.n1097 18.7549
R4612 VSS.n754 VSS.n748 18.4476
R4613 VSS.n1626 VSS.n888 18.4476
R4614 VSS.n864 VSS.t4 18.234
R4615 VSS.n1845 VSS.n844 18.0711
R4616 VSS.n1650 VSS.n1649 18.0711
R4617 VSS.t177 VSS.n1305 17.713
R4618 VSS.t178 VSS.n1629 17.713
R4619 VSS.t179 VSS.n782 17.713
R4620 VSS.n22 VSS.n10 17.3181
R4621 VSS.n982 VSS.n981 17.3181
R4622 VSS.n948 VSS.n924 17.3181
R4623 VSS.n719 VSS.n708 17.3181
R4624 VSS.n685 VSS.n684 17.3181
R4625 VSS.n975 VSS.n974 17.1928
R4626 VSS.n953 VSS.n920 17.1928
R4627 VSS.n712 VSS.n711 17.1928
R4628 VSS.n691 VSS.n690 17.1928
R4629 VSS.t2 VSS.n1543 17.1921
R4630 VSS.n1299 VSS.n1226 16.6711
R4631 VSS.n1322 VSS.n1232 16.6711
R4632 VSS.n1321 VSS.n1305 16.6711
R4633 VSS.n1310 VSS.n1309 16.6711
R4634 VSS.n1519 VSS.n1110 16.6711
R4635 VSS.n1530 VSS.n1106 16.6711
R4636 VSS.n1529 VSS.n1528 16.6711
R4637 VSS.n1537 VSS.n1536 16.6711
R4638 VSS.n1544 VSS.n1097 16.6711
R4639 VSS.n2106 VSS.n2105 16.6319
R4640 VSS.n29 VSS.n28 16.3559
R4641 VSS.n1299 VSS.t9 16.1502
R4642 VSS.n24 VSS.n11 15.8123
R4643 VSS.n978 VSS.n972 15.8123
R4644 VSS.n949 VSS.n922 15.8123
R4645 VSS.n716 VSS.n715 15.8123
R4646 VSS.n688 VSS.n659 15.8123
R4647 VSS.n1609 VSS.n1022 15.6292
R4648 VSS.n1616 VSS.n905 15.6292
R4649 VSS.n1637 VSS.n1636 15.6292
R4650 VSS.n907 VSS.n901 15.6292
R4651 VSS.n1629 VSS.n896 15.6292
R4652 VSS.n1655 VSS.n1654 15.6292
R4653 VSS.n1663 VSS.n890 15.6292
R4654 VSS.n1669 VSS.n885 15.6292
R4655 VSS.n1670 VSS.n868 15.6292
R4656 VSS.n2315 VSS.t54 15.1082
R4657 VSS.n2426 VSS.t84 15.1082
R4658 VSS.n1718 VSS.n1717 15.1082
R4659 VSS.n1016 VSS.n1015 15.0102
R4660 VSS.n368 VSS.n357 14.5711
R4661 VSS.n372 VSS.n371 14.5711
R4662 VSS.n355 VSS.n354 14.5711
R4663 VSS.n475 VSS.n474 14.5711
R4664 VSS.n471 VSS.n460 14.5711
R4665 VSS.n453 VSS.n452 14.5711
R4666 VSS.n427 VSS.n384 14.5711
R4667 VSS.n414 VSS.n330 14.5711
R4668 VSS.n113 VSS.n112 14.5711
R4669 VSS.n98 VSS.n92 14.5711
R4670 VSS.n72 VSS.n71 14.5711
R4671 VSS.n52 VSS.n44 14.5711
R4672 VSS.n977 VSS.n974 14.3064
R4673 VSS.n953 VSS.n952 14.3064
R4674 VSS.n712 VSS.n710 14.3064
R4675 VSS.n690 VSS.n689 14.3064
R4676 VSS.t42 VSS.n206 14.0663
R4677 VSS.n2378 VSS.t26 14.0663
R4678 VSS.n1844 VSS.n1842 13.5534
R4679 VSS.n1652 VSS.n1651 13.5534
R4680 VSS.n1601 VSS.t0 13.5454
R4681 VSS.n2108 VSS.n645 13.177
R4682 VSS.n2309 VSS.t16 13.0244
R4683 VSS.n166 VSS.t13 13.0244
R4684 VSS.n1740 VSS.t5 13.0244
R4685 VSS.n421 VSS.n333 12.7256
R4686 VSS.n419 VSS.n333 12.7256
R4687 VSS.n30 VSS.n4 12.7256
R4688 VSS.n1740 VSS.n857 12.5035
R4689 VSS.n1799 VSS.n1798 12.5035
R4690 VSS.n1798 VSS.t176 12.5035
R4691 VSS.n859 VSS.n852 12.5035
R4692 VSS.n1805 VSS.n853 12.5035
R4693 VSS.n1807 VSS.n825 12.5035
R4694 VSS.n1879 VSS.n1878 12.5035
R4695 VSS.n2109 VSS.n2108 12.424
R4696 VSS.n1845 VSS.n1844 12.0476
R4697 VSS.n1651 VSS.n1650 12.0476
R4698 VSS.n1591 VSS.n1080 11.9825
R4699 VSS.n1643 VSS.t7 11.9825
R4700 VSS.n12 VSS.n11 11.2946
R4701 VSS.n978 VSS.n977 11.2946
R4702 VSS.n952 VSS.n922 11.2946
R4703 VSS.n715 VSS.n710 11.2946
R4704 VSS.n689 VSS.n688 11.2946
R4705 VSS.n1003 VSS.n1002 11.0636
R4706 VSS.n1004 VSS.n962 11.0636
R4707 VSS.n1005 VSS.n961 11.0636
R4708 VSS.n1006 VSS.n914 11.0636
R4709 VSS.n955 VSS.n919 11.0636
R4710 VSS.n957 VSS.n956 11.0636
R4711 VSS.n959 VSS.n958 11.0636
R4712 VSS.n960 VSS.n913 11.0636
R4713 VSS.n1008 VSS.n1007 11.0636
R4714 VSS.n740 VSS.n739 11.0636
R4715 VSS.n741 VSS.n699 11.0636
R4716 VSS.n742 VSS.n698 11.0636
R4717 VSS.n743 VSS.n651 11.0636
R4718 VSS.n692 VSS.n656 11.0636
R4719 VSS.n694 VSS.n693 11.0636
R4720 VSS.n696 VSS.n695 11.0636
R4721 VSS.n697 VSS.n650 11.0636
R4722 VSS.n745 VSS.n744 11.0636
R4723 VSS.n1592 VSS.t0 10.9406
R4724 VSS.n1601 VSS.n1600 10.9406
R4725 VSS.t3 VSS.n1328 10.4196
R4726 VSS.n1528 VSS.t173 10.4196
R4727 VSS.t174 VSS.n1616 10.4196
R4728 VSS.t176 VSS.n859 10.4196
R4729 VSS.n1870 VSS.t91 10.4196
R4730 VSS.t1 VSS.n1106 9.89868
R4731 VSS.n1789 VSS.t5 9.89868
R4732 VSS.n24 VSS.n10 9.78874
R4733 VSS.n981 VSS.n972 9.78874
R4734 VSS.n949 VSS.n948 9.78874
R4735 VSS.n716 VSS.n708 9.78874
R4736 VSS.n685 VSS.n659 9.78874
R4737 VSS.n2549 VSS.n31 9.77955
R4738 VSS.n996 VSS.n964 9.58499
R4739 VSS.n933 VSS.n932 9.58499
R4740 VSS.n732 VSS.n700 9.58499
R4741 VSS.n669 VSS.n667 9.58499
R4742 VSS.n2107 VSS.n643 9.52595
R4743 VSS.n2502 VSS.n2501 9.49023
R4744 VSS.n327 VSS.n272 9.49023
R4745 VSS.n1626 VSS.n1625 9.49023
R4746 VSS.n1621 VSS.n1012 9.49023
R4747 VSS.n2102 VSS.n748 9.49023
R4748 VSS.n1493 VSS.n1484 9.49023
R4749 VSS.n1651 VSS.n1 9.36151
R4750 VSS.n1523 VSS.n2 9.36002
R4751 VSS.n1524 VSS.n2 9.36002
R4752 VSS.n1649 VSS.n1 9.35854
R4753 VSS.n359 VSS.n358 9.3005
R4754 VSS.n337 VSS.n336 9.3005
R4755 VSS.n351 VSS.n350 9.3005
R4756 VSS.n349 VSS.n348 9.3005
R4757 VSS.n343 VSS.n342 9.3005
R4758 VSS.n365 VSS.n364 9.3005
R4759 VSS.n367 VSS.n366 9.3005
R4760 VSS.n468 VSS.n467 9.3005
R4761 VSS.n470 VSS.n469 9.3005
R4762 VSS.n449 VSS.n448 9.3005
R4763 VSS.n447 VSS.n446 9.3005
R4764 VSS.n441 VSS.n440 9.3005
R4765 VSS.n463 VSS.n462 9.3005
R4766 VSS.n455 VSS.n454 9.3005
R4767 VSS.n422 VSS.n421 9.3005
R4768 VSS.n424 VSS.n423 9.3005
R4769 VSS.n426 VSS.n425 9.3005
R4770 VSS.n420 VSS.n419 9.3005
R4771 VSS.n418 VSS.n417 9.3005
R4772 VSS.n416 VSS.n415 9.3005
R4773 VSS.n4 VSS.n3 9.3005
R4774 VSS.n15 VSS.n14 9.3005
R4775 VSS.n17 VSS.n16 9.3005
R4776 VSS.n19 VSS.n18 9.3005
R4777 VSS.n21 VSS.n20 9.3005
R4778 VSS.n23 VSS.n22 9.3005
R4779 VSS.n25 VSS.n24 9.3005
R4780 VSS.n26 VSS.n12 9.3005
R4781 VSS.n95 VSS.n94 9.3005
R4782 VSS.n97 VSS.n96 9.3005
R4783 VSS.n107 VSS.n106 9.3005
R4784 VSS.n109 VSS.n108 9.3005
R4785 VSS.n86 VSS.n85 9.3005
R4786 VSS.n60 VSS.n50 9.3005
R4787 VSS.n53 VSS.n51 9.3005
R4788 VSS.n55 VSS.n54 9.3005
R4789 VSS.n68 VSS.n67 9.3005
R4790 VSS.n46 VSS.n45 9.3005
R4791 VSS.n480 VSS.n479 9.3005
R4792 VSS.n478 VSS.n269 9.3005
R4793 VSS.n327 VSS.n326 9.3005
R4794 VSS.n2497 VSS.n116 9.3005
R4795 VSS.n2501 VSS.n2500 9.3005
R4796 VSS.n2546 VSS.n2545 9.3005
R4797 VSS.n1843 VSS.n844 9.3005
R4798 VSS.n1844 VSS.n1843 9.3005
R4799 VSS.n964 VSS.n963 9.3005
R4800 VSS.n993 VSS.n992 9.3005
R4801 VSS.n991 VSS.n990 9.3005
R4802 VSS.n968 VSS.n967 9.3005
R4803 VSS.n985 VSS.n984 9.3005
R4804 VSS.n983 VSS.n982 9.3005
R4805 VSS.n972 VSS.n971 9.3005
R4806 VSS.n977 VSS.n976 9.3005
R4807 VSS.n934 VSS.n933 9.3005
R4808 VSS.n936 VSS.n935 9.3005
R4809 VSS.n928 VSS.n927 9.3005
R4810 VSS.n942 VSS.n941 9.3005
R4811 VSS.n944 VSS.n943 9.3005
R4812 VSS.n924 VSS.n923 9.3005
R4813 VSS.n950 VSS.n949 9.3005
R4814 VSS.n952 VSS.n951 9.3005
R4815 VSS.n733 VSS.n732 9.3005
R4816 VSS.n702 VSS.n701 9.3005
R4817 VSS.n727 VSS.n726 9.3005
R4818 VSS.n725 VSS.n724 9.3005
R4819 VSS.n706 VSS.n705 9.3005
R4820 VSS.n719 VSS.n718 9.3005
R4821 VSS.n717 VSS.n716 9.3005
R4822 VSS.n710 VSS.n709 9.3005
R4823 VSS.n667 VSS.n666 9.3005
R4824 VSS.n673 VSS.n672 9.3005
R4825 VSS.n675 VSS.n674 9.3005
R4826 VSS.n663 VSS.n662 9.3005
R4827 VSS.n681 VSS.n680 9.3005
R4828 VSS.n684 VSS.n683 9.3005
R4829 VSS.n682 VSS.n659 9.3005
R4830 VSS.n689 VSS.n658 9.3005
R4831 VSS.n1494 VSS.n1493 9.3005
R4832 VSS.n1485 VSS.n747 9.3005
R4833 VSS.n2102 VSS.n2101 9.3005
R4834 VSS.n1625 VSS.n1011 9.3005
R4835 VSS.n1634 VSS.n1010 9.3005
R4836 VSS.n1621 VSS.n1620 9.3005
R4837 VSS.n2106 VSS.n639 9.3005
R4838 VSS.n2108 VSS.n2107 9.3005
R4839 VSS.n1519 VSS.t1 8.85676
R4840 VSS.n399 VSS.n43 8.61608
R4841 VSS.n1537 VSS.t173 8.33581
R4842 VSS.n1024 VSS.n1015 8.33581
R4843 VSS.n22 VSS.n9 8.28285
R4844 VSS.n982 VSS.n970 8.28285
R4845 VSS.n945 VSS.n924 8.28285
R4846 VSS.n720 VSS.n719 8.28285
R4847 VSS.n684 VSS.n661 8.28285
R4848 VSS.n352 VSS.n347 8.2073
R4849 VSS.n450 VSS.n445 8.2073
R4850 VSS.n2328 VSS.t81 7.81485
R4851 VSS.n2414 VSS.t39 7.81485
R4852 VSS.n1788 VSS.n1787 7.81485
R4853 VSS.n844 VSS.n842 7.52991
R4854 VSS.n1649 VSS.n1648 7.52991
R4855 VSS.t111 VSS.n1016 7.50537
R4856 VSS.t7 VSS.n752 7.50537
R4857 VSS.n1617 VSS.n1015 7.29389
R4858 VSS.n1623 VSS.n646 7.25768
R4859 VSS.n2105 VSS.n2104 7.25768
R4860 VSS.n2100 VSS.n748 7.15344
R4861 VSS.n1627 VSS.n1626 7.15344
R4862 VSS.n20 VSS.n8 6.77697
R4863 VSS.n986 VSS.n985 6.77697
R4864 VSS.n944 VSS.n926 6.77697
R4865 VSS.n723 VSS.n706 6.77697
R4866 VSS.n680 VSS.n679 6.77697
R4867 VSS.t75 VSS.n214 6.77294
R4868 VSS.n2390 VSS.t63 6.77294
R4869 VSS.n363 VSS.n340 6.41949
R4870 VSS.n360 VSS.n338 6.41949
R4871 VSS.n464 VSS.n456 6.41949
R4872 VSS.n466 VSS.n458 6.41949
R4873 VSS.n93 VSS.n90 6.41949
R4874 VSS.n66 VSS.n47 6.41949
R4875 VSS.n1329 VSS.t3 6.25198
R4876 VSS.t158 VSS.n369 5.8005
R4877 VSS.n369 VSS.t60 5.8005
R4878 VSS.n370 VSS.t132 5.8005
R4879 VSS.n370 VSS.t158 5.8005
R4880 VSS.n353 VSS.t136 5.8005
R4881 VSS.n353 VSS.t32 5.8005
R4882 VSS.n473 VSS.t99 5.8005
R4883 VSS.n473 VSS.t97 5.8005
R4884 VSS.t97 VSS.n472 5.8005
R4885 VSS.n472 VSS.t17 5.8005
R4886 VSS.n451 VSS.t67 5.8005
R4887 VSS.n451 VSS.t70 5.8005
R4888 VSS.n374 VSS.t144 5.8005
R4889 VSS.n374 VSS.t14 5.8005
R4890 VSS.n378 VSS.t58 5.8005
R4891 VSS.n378 VSS.t120 5.8005
R4892 VSS.t27 VSS.n383 5.8005
R4893 VSS.n383 VSS.t64 5.8005
R4894 VSS.n429 VSS.t138 5.8005
R4895 VSS.n429 VSS.t170 5.8005
R4896 VSS.n433 VSS.t134 5.8005
R4897 VSS.n433 VSS.t142 5.8005
R4898 VSS.n437 VSS.t105 5.8005
R4899 VSS.n437 VSS.t55 5.8005
R4900 VSS.n376 VSS.t140 5.8005
R4901 VSS.n376 VSS.t168 5.8005
R4902 VSS.n380 VSS.t95 5.8005
R4903 VSS.n380 VSS.t89 5.8005
R4904 VSS.n328 VSS.t43 5.8005
R4905 VSS.n328 VSS.t50 5.8005
R4906 VSS.n431 VSS.t164 5.8005
R4907 VSS.n431 VSS.t162 5.8005
R4908 VSS.n435 VSS.t87 5.8005
R4909 VSS.n435 VSS.t160 5.8005
R4910 VSS.t170 VSS.n428 5.8005
R4911 VSS.n428 VSS.t27 5.8005
R4912 VSS.n99 VSS.t37 5.8005
R4913 VSS.t73 VSS.n99 5.8005
R4914 VSS.n100 VSS.t73 5.8005
R4915 VSS.n100 VSS.t127 5.8005
R4916 VSS.n82 VSS.t40 5.8005
R4917 VSS.n82 VSS.t85 5.8005
R4918 VSS.n80 VSS.t152 5.8005
R4919 VSS.n80 VSS.t150 5.8005
R4920 VSS.n78 VSS.t114 5.8005
R4921 VSS.n78 VSS.t125 5.8005
R4922 VSS.n76 VSS.t79 5.8005
R4923 VSS.n76 VSS.t76 5.8005
R4924 VSS.n74 VSS.t118 5.8005
R4925 VSS.n74 VSS.t82 5.8005
R4926 VSS.n70 VSS.t154 5.8005
R4927 VSS.n70 VSS.t35 5.8005
R4928 VSS.n63 VSS.t156 5.8005
R4929 VSS.n63 VSS.t154 5.8005
R4930 VSS.n2296 VSS.t69 5.73102
R4931 VSS.n158 VSS.t72 5.73102
R4932 VSS.t111 VSS.t174 5.73102
R4933 VSS.t6 VSS.t45 5.73102
R4934 VSS.n273 VSS.n272 5.64756
R4935 VSS.n2502 VSS.n2493 5.64756
R4936 VSS.n107 VSS.n103 5.37662
R4937 VSS.n62 VSS.n50 5.37662
R4938 VSS.n1471 VSS.t9 5.36112
R4939 VSS.n2072 VSS.t8 5.36112
R4940 VSS.n18 VSS.n7 5.27109
R4941 VSS.n989 VSS.n968 5.27109
R4942 VSS.n941 VSS.n940 5.27109
R4943 VSS.n724 VSS.n704 5.27109
R4944 VSS.n676 VSS.n663 5.27109
R4945 VSS.n886 VSS.t6 5.21007
R4946 VSS.n1879 VSS.t179 5.21007
R4947 VSS.n2290 VSS.n2289 4.68911
R4948 VSS.n1662 VSS.t45 4.68911
R4949 VSS.n1623 VSS.n1622 4.5683
R4950 VSS.n2104 VSS.n647 4.5683
R4951 VSS.n481 VSS.n480 4.51815
R4952 VSS.n2497 VSS.n117 4.51815
R4953 VSS.n1624 VSS.n1623 4.5005
R4954 VSS.n2104 VSS.n2103 4.5005
R4955 VSS.n2548 VSS.n114 4.26732
R4956 VSS.n1294 VSS.n1168 4.16815
R4957 VSS.n73 VSS.n44 3.81995
R4958 VSS.n367 VSS.n341 3.76521
R4959 VSS.n339 VSS.n337 3.76521
R4960 VSS.n344 VSS.n343 3.76521
R4961 VSS.n457 VSS.n455 3.76521
R4962 VSS.n470 VSS.n459 3.76521
R4963 VSS.n442 VSS.n441 3.76521
R4964 VSS.n426 VSS.n335 3.76521
R4965 VSS.n415 VSS.n331 3.76521
R4966 VSS.n16 VSS.n6 3.76521
R4967 VSS.n110 VSS.n86 3.76521
R4968 VSS.n97 VSS.n91 3.76521
R4969 VSS.n69 VSS.n46 3.76521
R4970 VSS.n56 VSS.n55 3.76521
R4971 VSS.n1526 VSS.n1523 3.76521
R4972 VSS.n990 VSS.n966 3.76521
R4973 VSS.n937 VSS.n928 3.76521
R4974 VSS.n728 VSS.n727 3.76521
R4975 VSS.n675 VSS.n665 3.76521
R4976 VSS.n2550 VSS.n2549 3.74842
R4977 VSS.n1617 VSS.t111 3.6472
R4978 VSS.n1630 VSS.t7 3.6472
R4979 VSS.n1495 VSS.n1494 3.38874
R4980 VSS.n1620 VSS.n1619 3.38874
R4981 VSS.n478 VSS.n477 3.11834
R4982 VSS.n976 VSS.n975 3.09986
R4983 VSS.n951 VSS.n920 3.09986
R4984 VSS.n711 VSS.n709 3.09986
R4985 VSS.n691 VSS.n658 3.09986
R4986 VSS.n1496 VSS.n1484 3.01226
R4987 VSS.n1013 VSS.n1012 3.01226
R4988 VSS.n373 VSS.n372 2.89851
R4989 VSS.n460 VSS.n439 2.89851
R4990 VSS VSS.n2551 2.69823
R4991 VSS.n92 VSS.n84 2.67025
R4992 VSS.n114 VSS.n113 2.67025
R4993 VSS.n73 VSS.n72 2.67025
R4994 VSS.n1232 VSS.t9 2.60528
R4995 VSS.n853 VSS.t8 2.60528
R4996 VSS.n2105 VSS.n646 2.5952
R4997 VSS.n29 VSS.t180 2.48621
R4998 VSS.n29 VSS.t92 2.48621
R4999 VSS.t146 VSS.n1003 2.48621
R5000 VSS.n1003 VSS.t23 2.48621
R5001 VSS.t103 VSS.n1004 2.48621
R5002 VSS.n1004 VSS.t146 2.48621
R5003 VSS.t48 VSS.n1005 2.48621
R5004 VSS.n1005 VSS.t103 2.48621
R5005 VSS.t109 VSS.n1006 2.48621
R5006 VSS.n1006 VSS.t48 2.48621
R5007 VSS.n955 VSS.t29 2.48621
R5008 VSS.t21 VSS.n955 2.48621
R5009 VSS.n956 VSS.t21 2.48621
R5010 VSS.n956 VSS.t11 2.48621
R5011 VSS.n959 VSS.t11 2.48621
R5012 VSS.t172 VSS.n959 2.48621
R5013 VSS.n960 VSS.t172 2.48621
R5014 VSS.t112 VSS.n960 2.48621
R5015 VSS.n1007 VSS.t112 2.48621
R5016 VSS.n1007 VSS.t109 2.48621
R5017 VSS.t116 VSS.n740 2.48621
R5018 VSS.n740 VSS.t122 2.48621
R5019 VSS.t101 VSS.n741 2.48621
R5020 VSS.n741 VSS.t116 2.48621
R5021 VSS.t46 VSS.n742 2.48621
R5022 VSS.n742 VSS.t101 2.48621
R5023 VSS.t166 VSS.n743 2.48621
R5024 VSS.n743 VSS.t46 2.48621
R5025 VSS.n692 VSS.t19 2.48621
R5026 VSS.t52 VSS.n692 2.48621
R5027 VSS.n693 VSS.t52 2.48621
R5028 VSS.n693 VSS.t107 2.48621
R5029 VSS.n696 VSS.t107 2.48621
R5030 VSS.t148 VSS.n696 2.48621
R5031 VSS.n697 VSS.t148 2.48621
R5032 VSS.t130 VSS.n697 2.48621
R5033 VSS.n744 VSS.t130 2.48621
R5034 VSS.n744 VSS.t166 2.48621
R5035 VSS.n28 VSS.n27 2.36936
R5036 VSS.n2547 VSS.n2546 2.33344
R5037 VSS.n348 VSS.n345 2.25932
R5038 VSS.n446 VSS.n443 2.25932
R5039 VSS.n423 VSS.n334 2.25932
R5040 VSS.n417 VSS.n332 2.25932
R5041 VSS.n14 VSS.n5 2.25932
R5042 VSS.n109 VSS.n88 2.25932
R5043 VSS.n59 VSS.n51 2.25932
R5044 VSS.n994 VSS.n993 2.25932
R5045 VSS.n936 VSS.n930 2.25932
R5046 VSS.n731 VSS.n702 2.25932
R5047 VSS.n672 VSS.n671 2.25932
R5048 VSS.n356 VSS.n115 2.25177
R5049 VSS.n477 VSS.n476 2.25177
R5050 VSS.n401 VSS.n400 2.25162
R5051 VSS.n403 VSS.n402 2.25162
R5052 VSS.n405 VSS.n404 2.25162
R5053 VSS.n407 VSS.n406 2.25162
R5054 VSS.n409 VSS.n408 2.25162
R5055 VSS.n398 VSS.n397 2.25162
R5056 VSS.n411 VSS.n410 2.25162
R5057 VSS.n395 VSS.n394 2.25162
R5058 VSS.n393 VSS.n392 2.25162
R5059 VSS.n391 VSS.n390 2.25162
R5060 VSS.n389 VSS.n388 2.25162
R5061 VSS.n387 VSS.n386 2.25162
R5062 VSS.n43 VSS.n42 2.17137
R5063 VSS.n1630 VSS.t178 2.08433
R5064 VSS.n1717 VSS.t4 2.08433
R5065 VSS.n2549 VSS.n43 1.94432
R5066 VSS.n2551 VSS.n2550 1.74238
R5067 VSS.n521 VSS.t66 1.56337
R5068 VSS.t31 VSS.n145 1.56337
R5069 VSS.n1544 VSS.t2 1.56337
R5070 VSS.n2549 VSS.n2548 1.33979
R5071 VSS.n75 VSS.n73 1.1502
R5072 VSS.n77 VSS.n75 1.1502
R5073 VSS.n79 VSS.n77 1.1502
R5074 VSS.n81 VSS.n79 1.1502
R5075 VSS.n83 VSS.n81 1.1502
R5076 VSS.n84 VSS.n83 1.1502
R5077 VSS.n114 VSS.n84 1.1502
R5078 VSS.n1310 VSS.t177 1.04241
R5079 VSS.n2548 VSS.n2547 0.805174
R5080 VSS.n2547 VSS.n115 0.7864
R5081 VSS.n1002 VSS.n997 0.779912
R5082 VSS.n1002 VSS.n962 0.779912
R5083 VSS.n962 VSS.n961 0.779912
R5084 VSS.n961 VSS.n914 0.779912
R5085 VSS.n931 VSS.n919 0.779912
R5086 VSS.n957 VSS.n919 0.779912
R5087 VSS.n958 VSS.n957 0.779912
R5088 VSS.n958 VSS.n913 0.779912
R5089 VSS.n1008 VSS.n913 0.779912
R5090 VSS.n1008 VSS.n914 0.779912
R5091 VSS.n739 VSS.n734 0.779912
R5092 VSS.n739 VSS.n699 0.779912
R5093 VSS.n699 VSS.n698 0.779912
R5094 VSS.n698 VSS.n651 0.779912
R5095 VSS.n668 VSS.n656 0.779912
R5096 VSS.n694 VSS.n656 0.779912
R5097 VSS.n695 VSS.n694 0.779912
R5098 VSS.n695 VSS.n650 0.779912
R5099 VSS.n745 VSS.n650 0.779912
R5100 VSS.n745 VSS.n651 0.779912
R5101 VSS.n106 VSS.n105 0.753441
R5102 VSS.n61 VSS.n60 0.753441
R5103 VSS.n326 VSS.n325 0.753441
R5104 VSS.n2500 VSS.n2496 0.753441
R5105 VSS.n1525 VSS.n1524 0.753441
R5106 VSS.n2101 VSS.n749 0.753441
R5107 VSS.n1632 VSS.n1011 0.753441
R5108 VSS.n998 VSS.n911 0.701719
R5109 VSS.n999 VSS.n998 0.701719
R5110 VSS.n1000 VSS.n999 0.701719
R5111 VSS.n917 VSS.n916 0.701719
R5112 VSS.n916 VSS.n915 0.701719
R5113 VSS.n915 VSS.n912 0.701719
R5114 VSS.n735 VSS.n648 0.701719
R5115 VSS.n736 VSS.n735 0.701719
R5116 VSS.n737 VSS.n736 0.701719
R5117 VSS.n654 VSS.n653 0.701719
R5118 VSS.n653 VSS.n652 0.701719
R5119 VSS.n652 VSS.n649 0.701719
R5120 VSS.n646 VSS.n0 0.675121
R5121 VSS.n357 VSS.n356 0.647239
R5122 VSS.n476 VSS.n475 0.647239
R5123 VSS.n389 VSS.n387 0.574917
R5124 VSS.n391 VSS.n389 0.574917
R5125 VSS.n393 VSS.n391 0.574917
R5126 VSS.n395 VSS.n393 0.574917
R5127 VSS.n398 VSS.n395 0.574917
R5128 VSS.n410 VSS.n398 0.574917
R5129 VSS.n410 VSS.n409 0.574917
R5130 VSS.n409 VSS.n407 0.574917
R5131 VSS.n407 VSS.n405 0.574917
R5132 VSS.n405 VSS.n403 0.574917
R5133 VSS.n403 VSS.n401 0.574917
R5134 VSS.n401 VSS.n399 0.574917
R5135 VSS.n33 VSS.n32 0.574917
R5136 VSS.n34 VSS.n33 0.574917
R5137 VSS.n35 VSS.n34 0.574917
R5138 VSS.n36 VSS.n35 0.574917
R5139 VSS.n37 VSS.n36 0.574917
R5140 VSS.n38 VSS.n37 0.574917
R5141 VSS.n39 VSS.n38 0.574917
R5142 VSS.n40 VSS.n39 0.574917
R5143 VSS.n41 VSS.n40 0.574917
R5144 VSS.n42 VSS.n41 0.574917
R5145 VSS.n477 VSS.n439 0.574311
R5146 VSS.n439 VSS.n438 0.574311
R5147 VSS.n438 VSS.n436 0.574311
R5148 VSS.n436 VSS.n434 0.574311
R5149 VSS.n434 VSS.n432 0.574311
R5150 VSS.n432 VSS.n430 0.574311
R5151 VSS.n430 VSS.n329 0.574311
R5152 VSS.n382 VSS.n329 0.574311
R5153 VSS.n382 VSS.n381 0.574311
R5154 VSS.n381 VSS.n379 0.574311
R5155 VSS.n379 VSS.n377 0.574311
R5156 VSS.n377 VSS.n375 0.574311
R5157 VSS.n375 VSS.n373 0.574311
R5158 VSS.n373 VSS.n115 0.574311
R5159 VSS.n2341 VSS.t78 0.521457
R5160 VSS.n2402 VSS.t57 0.521457
R5161 VSS.n356 VSS.n355 0.418978
R5162 VSS.n476 VSS.n453 0.418978
R5163 VSS.n1001 VSS.n1000 0.35111
R5164 VSS.n918 VSS.n917 0.35111
R5165 VSS.n738 VSS.n737 0.35111
R5166 VSS.n655 VSS.n654 0.35111
R5167 VSS VSS.n0 0.3505
R5168 VSS.n361 VSS.n360 0.320353
R5169 VSS.n363 VSS.n361 0.320353
R5170 VSS.n363 VSS.n362 0.320353
R5171 VSS.n347 VSS.n346 0.320353
R5172 VSS.n466 VSS.n465 0.320353
R5173 VSS.n464 VSS.n461 0.320353
R5174 VSS.n465 VSS.n464 0.320353
R5175 VSS.n445 VSS.n444 0.320353
R5176 VSS.n27 VSS.n13 0.320353
R5177 VSS.n93 VSS.n89 0.320353
R5178 VSS.n101 VSS.n89 0.320353
R5179 VSS.n102 VSS.n101 0.320353
R5180 VSS.n107 VSS.n102 0.320353
R5181 VSS.n50 VSS.n48 0.320353
R5182 VSS.n64 VSS.n48 0.320353
R5183 VSS.n65 VSS.n64 0.320353
R5184 VSS.n66 VSS.n65 0.320353
R5185 VSS.n2550 VSS.n2 0.303278
R5186 VSS.n2551 VSS.n1 0.303278
R5187 VSS.n396 VSS.n385 0.302413
R5188 VSS.n412 VSS.n385 0.302413
R5189 VSS.n1009 VSS.n1008 0.272321
R5190 VSS.n746 VSS.n745 0.272321
R5191 VSS.n1009 VSS.n911 0.261436
R5192 VSS.n1009 VSS.n912 0.261436
R5193 VSS.n746 VSS.n648 0.261436
R5194 VSS.n746 VSS.n649 0.261436
R5195 VSS.n1002 VSS.n1001 0.228761
R5196 VSS.n919 VSS.n918 0.228761
R5197 VSS.n739 VSS.n738 0.228761
R5198 VSS.n656 VSS.n655 0.228761
R5199 VSS.n2107 VSS.n2106 0.21925
R5200 VSS.n385 VSS.n384 0.217891
R5201 VSS.n414 VSS.n413 0.217891
R5202 VSS.n1625 VSS.n1624 0.217762
R5203 VSS.n2103 VSS.n2102 0.217762
R5204 VSS.n2501 VSS.n116 0.204927
R5205 VSS.n479 VSS.n327 0.204927
R5206 VSS.n372 VSS.n336 0.196152
R5207 VSS.n359 VSS.n336 0.196152
R5208 VSS.n360 VSS.n359 0.196152
R5209 VSS.n350 VSS.n347 0.196152
R5210 VSS.n350 VSS.n349 0.196152
R5211 VSS.n349 VSS.n342 0.196152
R5212 VSS.n355 VSS.n342 0.196152
R5213 VSS.n366 VSS.n357 0.196152
R5214 VSS.n366 VSS.n365 0.196152
R5215 VSS.n365 VSS.n363 0.196152
R5216 VSS.n469 VSS.n460 0.196152
R5217 VSS.n469 VSS.n468 0.196152
R5218 VSS.n468 VSS.n466 0.196152
R5219 VSS.n448 VSS.n445 0.196152
R5220 VSS.n448 VSS.n447 0.196152
R5221 VSS.n447 VSS.n440 0.196152
R5222 VSS.n453 VSS.n440 0.196152
R5223 VSS.n475 VSS.n454 0.196152
R5224 VSS.n463 VSS.n454 0.196152
R5225 VSS.n464 VSS.n463 0.196152
R5226 VSS.n425 VSS.n384 0.196152
R5227 VSS.n425 VSS.n424 0.196152
R5228 VSS.n424 VSS.n422 0.196152
R5229 VSS.n422 VSS.n420 0.196152
R5230 VSS.n420 VSS.n418 0.196152
R5231 VSS.n418 VSS.n416 0.196152
R5232 VSS.n416 VSS.n414 0.196152
R5233 VSS.n27 VSS.n26 0.196152
R5234 VSS.n26 VSS.n25 0.196152
R5235 VSS.n25 VSS.n23 0.196152
R5236 VSS.n23 VSS.n21 0.196152
R5237 VSS.n21 VSS.n19 0.196152
R5238 VSS.n19 VSS.n17 0.196152
R5239 VSS.n17 VSS.n15 0.196152
R5240 VSS.n15 VSS.n3 0.196152
R5241 VSS.n31 VSS.n3 0.196152
R5242 VSS.n96 VSS.n92 0.196152
R5243 VSS.n96 VSS.n95 0.196152
R5244 VSS.n95 VSS.n93 0.196152
R5245 VSS.n113 VSS.n85 0.196152
R5246 VSS.n108 VSS.n85 0.196152
R5247 VSS.n108 VSS.n107 0.196152
R5248 VSS.n54 VSS.n44 0.196152
R5249 VSS.n54 VSS.n53 0.196152
R5250 VSS.n53 VSS.n50 0.196152
R5251 VSS.n72 VSS.n45 0.196152
R5252 VSS.n67 VSS.n45 0.196152
R5253 VSS.n67 VSS.n66 0.196152
R5254 VSS.n976 VSS.n971 0.196152
R5255 VSS.n983 VSS.n971 0.196152
R5256 VSS.n984 VSS.n983 0.196152
R5257 VSS.n984 VSS.n967 0.196152
R5258 VSS.n991 VSS.n967 0.196152
R5259 VSS.n992 VSS.n991 0.196152
R5260 VSS.n992 VSS.n963 0.196152
R5261 VSS.n997 VSS.n963 0.196152
R5262 VSS.n951 VSS.n950 0.196152
R5263 VSS.n950 VSS.n923 0.196152
R5264 VSS.n943 VSS.n923 0.196152
R5265 VSS.n943 VSS.n942 0.196152
R5266 VSS.n942 VSS.n927 0.196152
R5267 VSS.n935 VSS.n927 0.196152
R5268 VSS.n935 VSS.n934 0.196152
R5269 VSS.n934 VSS.n931 0.196152
R5270 VSS.n734 VSS.n733 0.196152
R5271 VSS.n733 VSS.n701 0.196152
R5272 VSS.n726 VSS.n701 0.196152
R5273 VSS.n726 VSS.n725 0.196152
R5274 VSS.n725 VSS.n705 0.196152
R5275 VSS.n718 VSS.n705 0.196152
R5276 VSS.n718 VSS.n717 0.196152
R5277 VSS.n717 VSS.n709 0.196152
R5278 VSS.n668 VSS.n666 0.196152
R5279 VSS.n673 VSS.n666 0.196152
R5280 VSS.n674 VSS.n673 0.196152
R5281 VSS.n674 VSS.n662 0.196152
R5282 VSS.n681 VSS.n662 0.196152
R5283 VSS.n683 VSS.n681 0.196152
R5284 VSS.n683 VSS.n682 0.196152
R5285 VSS.n682 VSS.n658 0.196152
R5286 VSS.n1622 VSS.n1621 0.193208
R5287 VSS.n1493 VSS.n647 0.193208
R5288 VSS.n397 VSS.n396 0.142018
R5289 VSS.n412 VSS.n411 0.142018
R5290 VSS.n1010 VSS.n1009 0.114136
R5291 VSS.n747 VSS.n746 0.114136
R5292 VSS.n2546 VSS.n116 0.104667
R5293 VSS.n479 VSS.n478 0.104667
R5294 VSS.n1843 VSS.n0 0.0771129
R5295 VSS.n1622 VSS.n1010 0.048119
R5296 VSS.n1624 VSS.n1010 0.048119
R5297 VSS.n747 VSS.n647 0.048119
R5298 VSS.n2103 VSS.n747 0.048119
R5299 a_4920_2896.n51 a_4920_2896.n6 185
R5300 a_4920_2896.n51 a_4920_2896.n4 185
R5301 a_4920_2896.n51 a_4920_2896.n7 185
R5302 a_4920_2896.n51 a_4920_2896.n3 185
R5303 a_4920_2896.n51 a_4920_2896.n8 185
R5304 a_4920_2896.n51 a_4920_2896.n2 185
R5305 a_4920_2896.n51 a_4920_2896.n50 185
R5306 a_4920_2896.n0 a_4920_2896.t0 130.75
R5307 a_4920_2896.t1 a_4920_2896.n0 91.3557
R5308 a_4920_2896.n51 a_4920_2896.n1 86.5152
R5309 a_4920_2896.n11 a_4920_2896.n5 30.3012
R5310 a_4920_2896.n30 a_4920_2896.n29 26.8581
R5311 a_4920_2896.n41 a_4920_2896.n40 26.6299
R5312 a_4920_2896.n34 a_4920_2896.n24 25.7063
R5313 a_4920_2896.n33 a_4920_2896.n25 25.7063
R5314 a_4920_2896.n32 a_4920_2896.n26 25.7063
R5315 a_4920_2896.n31 a_4920_2896.n27 25.7063
R5316 a_4920_2896.n30 a_4920_2896.n28 25.7063
R5317 a_4920_2896.n41 a_4920_2896.n39 25.4781
R5318 a_4920_2896.n42 a_4920_2896.n38 25.4781
R5319 a_4920_2896.n43 a_4920_2896.n37 25.4781
R5320 a_4920_2896.n44 a_4920_2896.n36 25.4781
R5321 a_4920_2896.n45 a_4920_2896.n35 25.4781
R5322 a_4920_2896.n50 a_4920_2896.n49 24.8476
R5323 a_4920_2896.n9 a_4920_2896.n2 23.3417
R5324 a_4920_2896.n47 a_4920_2896.n1 22.0256
R5325 a_4920_2896.n21 a_4920_2896.n8 21.8358
R5326 a_4920_2896.n19 a_4920_2896.n3 20.3299
R5327 a_4920_2896.n17 a_4920_2896.n7 18.824
R5328 a_4920_2896.n15 a_4920_2896.n4 17.3181
R5329 a_4920_2896.n51 a_4920_2896.n5 16.3559
R5330 a_4920_2896.n13 a_4920_2896.n6 15.8123
R5331 a_4920_2896.n49 a_4920_2896.n1 12.7256
R5332 a_4920_2896.n11 a_4920_2896.n6 11.2946
R5333 a_4920_2896.n13 a_4920_2896.n4 9.78874
R5334 a_4920_2896.n46 a_4920_2896.n34 9.30285
R5335 a_4920_2896.n49 a_4920_2896.n48 9.3005
R5336 a_4920_2896.n23 a_4920_2896.n9 9.3005
R5337 a_4920_2896.n22 a_4920_2896.n21 9.3005
R5338 a_4920_2896.n20 a_4920_2896.n19 9.3005
R5339 a_4920_2896.n18 a_4920_2896.n17 9.3005
R5340 a_4920_2896.n16 a_4920_2896.n15 9.3005
R5341 a_4920_2896.n14 a_4920_2896.n13 9.3005
R5342 a_4920_2896.n12 a_4920_2896.n11 9.3005
R5343 a_4920_2896.n15 a_4920_2896.n7 8.28285
R5344 a_4920_2896.n17 a_4920_2896.n3 6.77697
R5345 a_4920_2896.n40 a_4920_2896.t16 5.8005
R5346 a_4920_2896.n40 a_4920_2896.t11 5.8005
R5347 a_4920_2896.n39 a_4920_2896.t24 5.8005
R5348 a_4920_2896.n39 a_4920_2896.t23 5.8005
R5349 a_4920_2896.n38 a_4920_2896.t22 5.8005
R5350 a_4920_2896.n38 a_4920_2896.t5 5.8005
R5351 a_4920_2896.n37 a_4920_2896.t6 5.8005
R5352 a_4920_2896.n37 a_4920_2896.t13 5.8005
R5353 a_4920_2896.n36 a_4920_2896.t12 5.8005
R5354 a_4920_2896.n36 a_4920_2896.t18 5.8005
R5355 a_4920_2896.n35 a_4920_2896.t25 5.8005
R5356 a_4920_2896.n35 a_4920_2896.t17 5.8005
R5357 a_4920_2896.n24 a_4920_2896.t10 5.8005
R5358 a_4920_2896.n24 a_4920_2896.t3 5.8005
R5359 a_4920_2896.n25 a_4920_2896.t20 5.8005
R5360 a_4920_2896.n25 a_4920_2896.t4 5.8005
R5361 a_4920_2896.n26 a_4920_2896.t15 5.8005
R5362 a_4920_2896.n26 a_4920_2896.t21 5.8005
R5363 a_4920_2896.n27 a_4920_2896.t7 5.8005
R5364 a_4920_2896.n27 a_4920_2896.t14 5.8005
R5365 a_4920_2896.n28 a_4920_2896.t9 5.8005
R5366 a_4920_2896.n28 a_4920_2896.t8 5.8005
R5367 a_4920_2896.n29 a_4920_2896.t2 5.8005
R5368 a_4920_2896.n29 a_4920_2896.t19 5.8005
R5369 a_4920_2896.n19 a_4920_2896.n8 5.27109
R5370 a_4920_2896.n21 a_4920_2896.n2 3.76521
R5371 a_4920_2896.n46 a_4920_2896.n45 2.92217
R5372 a_4920_2896.t1 a_4920_2896.n51 2.48621
R5373 a_4920_2896.n51 a_4920_2896.t26 2.48621
R5374 a_4920_2896.n10 a_4920_2896.n5 2.36936
R5375 a_4920_2896.n50 a_4920_2896.n9 2.25932
R5376 a_4920_2896.n47 a_4920_2896.n46 2.19829
R5377 a_4920_2896.n42 a_4920_2896.n41 1.15229
R5378 a_4920_2896.n43 a_4920_2896.n42 1.15229
R5379 a_4920_2896.n44 a_4920_2896.n43 1.15229
R5380 a_4920_2896.n45 a_4920_2896.n44 1.15229
R5381 a_4920_2896.n31 a_4920_2896.n30 1.15229
R5382 a_4920_2896.n32 a_4920_2896.n31 1.15229
R5383 a_4920_2896.n33 a_4920_2896.n32 1.15229
R5384 a_4920_2896.n34 a_4920_2896.n33 1.15229
R5385 a_4920_2896.n10 a_4920_2896.n0 0.320353
R5386 a_4920_2896.n12 a_4920_2896.n10 0.196152
R5387 a_4920_2896.n14 a_4920_2896.n12 0.196152
R5388 a_4920_2896.n16 a_4920_2896.n14 0.196152
R5389 a_4920_2896.n18 a_4920_2896.n16 0.196152
R5390 a_4920_2896.n20 a_4920_2896.n18 0.196152
R5391 a_4920_2896.n22 a_4920_2896.n20 0.196152
R5392 a_4920_2896.n23 a_4920_2896.n22 0.196152
R5393 a_4920_2896.n48 a_4920_2896.n23 0.196152
R5394 a_4920_2896.n48 a_4920_2896.n47 0.196152
R5395 VP.n0 VP.t7 263.647
R5396 VP.n3 VP.t3 262.863
R5397 VP.n2 VP.t1 262.498
R5398 VP.n0 VP.t6 261.709
R5399 VP.n1 VP.t2 261.709
R5400 VP.n3 VP.t5 261.584
R5401 VP.n4 VP.t4 261.584
R5402 VP.n5 VP.t0 261.433
R5403 VP.n6 VP.n2 8.91142
R5404 VP VP.n6 2.39915
R5405 VP.n1 VP.n0 1.72698
R5406 VP.n6 VP.n5 1.52193
R5407 VP.n5 VP.n4 1.4312
R5408 VP.n4 VP.n3 1.16675
R5409 VP.n2 VP.n1 1.14999
R5410 a_2995_7336.n32 a_2995_7336.n31 185
R5411 a_2995_7336.n32 a_2995_7336.n14 185
R5412 a_2995_7336.n32 a_2995_7336.n13 185
R5413 a_2995_7336.n32 a_2995_7336.n12 185
R5414 a_2995_7336.n32 a_2995_7336.n11 185
R5415 a_2995_7336.n32 a_2995_7336.n10 185
R5416 a_2995_7336.n32 a_2995_7336.n9 185
R5417 a_2995_7336.n15 a_2995_7336.t9 130.75
R5418 a_2995_7336.n15 a_2995_7336.t11 91.3557
R5419 a_2995_7336.n33 a_2995_7336.n32 86.5152
R5420 a_2995_7336.n17 a_2995_7336.n8 30.3012
R5421 a_2995_7336.n31 a_2995_7336.n7 24.8476
R5422 a_2995_7336.n30 a_2995_7336.n14 23.3417
R5423 a_2995_7336.n34 a_2995_7336.n33 22.0256
R5424 a_2995_7336.n27 a_2995_7336.n13 21.8358
R5425 a_2995_7336.n25 a_2995_7336.n12 20.3299
R5426 a_2995_7336.n23 a_2995_7336.n11 18.824
R5427 a_2995_7336.n21 a_2995_7336.n10 17.3181
R5428 a_2995_7336.n32 a_2995_7336.n8 16.3559
R5429 a_2995_7336.n19 a_2995_7336.n9 15.8123
R5430 a_2995_7336.n33 a_2995_7336.n7 12.7256
R5431 a_2995_7336.n38 a_2995_7336.n37 12.1709
R5432 a_2995_7336.n39 a_2995_7336.n38 12.1709
R5433 a_2995_7336.n41 a_2995_7336.n40 11.4939
R5434 a_2995_7336.n37 a_2995_7336.n35 11.493
R5435 a_2995_7336.n3 a_2995_7336.n1 11.493
R5436 a_2995_7336.n39 a_2995_7336.n4 11.493
R5437 a_2995_7336.n40 a_2995_7336.n0 11.4929
R5438 a_2995_7336.n37 a_2995_7336.n36 11.4929
R5439 a_2995_7336.n3 a_2995_7336.n2 11.4929
R5440 a_2995_7336.n39 a_2995_7336.n5 11.4929
R5441 a_2995_7336.n17 a_2995_7336.n9 11.2946
R5442 a_2995_7336.n19 a_2995_7336.n10 9.78874
R5443 a_2995_7336.n7 a_2995_7336.n6 9.3005
R5444 a_2995_7336.n30 a_2995_7336.n29 9.3005
R5445 a_2995_7336.n28 a_2995_7336.n27 9.3005
R5446 a_2995_7336.n26 a_2995_7336.n25 9.3005
R5447 a_2995_7336.n24 a_2995_7336.n23 9.3005
R5448 a_2995_7336.n22 a_2995_7336.n21 9.3005
R5449 a_2995_7336.n20 a_2995_7336.n19 9.3005
R5450 a_2995_7336.n18 a_2995_7336.n17 9.3005
R5451 a_2995_7336.n21 a_2995_7336.n11 8.28285
R5452 a_2995_7336.n23 a_2995_7336.n12 6.77697
R5453 a_2995_7336.n25 a_2995_7336.n13 5.27109
R5454 a_2995_7336.n27 a_2995_7336.n14 3.76521
R5455 a_2995_7336.n38 a_2995_7336.n34 3.48602
R5456 a_2995_7336.n0 a_2995_7336.t3 2.48621
R5457 a_2995_7336.n0 a_2995_7336.t18 2.48621
R5458 a_2995_7336.n36 a_2995_7336.t8 2.48621
R5459 a_2995_7336.n36 a_2995_7336.t14 2.48621
R5460 a_2995_7336.n35 a_2995_7336.t15 2.48621
R5461 a_2995_7336.n35 a_2995_7336.t7 2.48621
R5462 a_2995_7336.n2 a_2995_7336.t19 2.48621
R5463 a_2995_7336.n2 a_2995_7336.t4 2.48621
R5464 a_2995_7336.n1 a_2995_7336.t6 2.48621
R5465 a_2995_7336.n1 a_2995_7336.t12 2.48621
R5466 a_2995_7336.n5 a_2995_7336.t13 2.48621
R5467 a_2995_7336.n5 a_2995_7336.t5 2.48621
R5468 a_2995_7336.n4 a_2995_7336.t1 2.48621
R5469 a_2995_7336.n4 a_2995_7336.t17 2.48621
R5470 a_2995_7336.n32 a_2995_7336.t16 2.48621
R5471 a_2995_7336.n32 a_2995_7336.t10 2.48621
R5472 a_2995_7336.t0 a_2995_7336.n41 2.48621
R5473 a_2995_7336.n41 a_2995_7336.t2 2.48621
R5474 a_2995_7336.n16 a_2995_7336.n8 2.36936
R5475 a_2995_7336.n31 a_2995_7336.n30 2.25932
R5476 a_2995_7336.n37 a_2995_7336.n3 1.15229
R5477 a_2995_7336.n40 a_2995_7336.n3 1.15229
R5478 a_2995_7336.n40 a_2995_7336.n39 1.15229
R5479 a_2995_7336.n16 a_2995_7336.n15 0.320353
R5480 a_2995_7336.n34 a_2995_7336.n6 0.196152
R5481 a_2995_7336.n29 a_2995_7336.n6 0.196152
R5482 a_2995_7336.n29 a_2995_7336.n28 0.196152
R5483 a_2995_7336.n28 a_2995_7336.n26 0.196152
R5484 a_2995_7336.n26 a_2995_7336.n24 0.196152
R5485 a_2995_7336.n24 a_2995_7336.n22 0.196152
R5486 a_2995_7336.n22 a_2995_7336.n20 0.196152
R5487 a_2995_7336.n20 a_2995_7336.n18 0.196152
R5488 a_2995_7336.n18 a_2995_7336.n16 0.196152
R5489 VN.n0 VN.t0 263.647
R5490 VN.n3 VN.t2 262.863
R5491 VN.n2 VN.t5 262.498
R5492 VN.n1 VN.t4 261.709
R5493 VN.n0 VN.t1 261.709
R5494 VN.n4 VN.t7 261.584
R5495 VN.n3 VN.t6 261.584
R5496 VN.n5 VN.t3 261.433
R5497 VN.n6 VN.n2 8.91142
R5498 VN VN.n6 2.48969
R5499 VN.n1 VN.n0 1.72698
R5500 VN.n6 VN.n5 1.52193
R5501 VN.n5 VN.n4 1.4312
R5502 VN.n4 VN.n3 1.16675
R5503 VN.n2 VN.n1 1.14999
R5504 a_2479_9004.n17 a_2479_9004.t22 260.111
R5505 a_2479_9004.n15 a_2479_9004.t21 260.111
R5506 a_2479_9004.n14 a_2479_9004.t5 260.111
R5507 a_2479_9004.n12 a_2479_9004.t7 260.111
R5508 a_2479_9004.n17 a_2479_9004.t9 260.111
R5509 a_2479_9004.n15 a_2479_9004.t11 260.111
R5510 a_2479_9004.n14 a_2479_9004.t24 260.111
R5511 a_2479_9004.n12 a_2479_9004.t23 260.111
R5512 a_2479_9004.n13 a_2479_9004.n11 203.413
R5513 a_2479_9004.n16 a_2479_9004.n10 203.413
R5514 a_2479_9004.n48 a_2479_9004.n47 185
R5515 a_2479_9004.n48 a_2479_9004.n30 185
R5516 a_2479_9004.n48 a_2479_9004.n29 185
R5517 a_2479_9004.n48 a_2479_9004.n28 185
R5518 a_2479_9004.n48 a_2479_9004.n27 185
R5519 a_2479_9004.n48 a_2479_9004.n26 185
R5520 a_2479_9004.n48 a_2479_9004.n25 185
R5521 a_2479_9004.n72 a_2479_9004.n4 185
R5522 a_2479_9004.n72 a_2479_9004.n6 185
R5523 a_2479_9004.n72 a_2479_9004.n3 185
R5524 a_2479_9004.n72 a_2479_9004.n7 185
R5525 a_2479_9004.n72 a_2479_9004.n2 185
R5526 a_2479_9004.n72 a_2479_9004.n8 185
R5527 a_2479_9004.n72 a_2479_9004.n1 185
R5528 a_2479_9004.n0 a_2479_9004.t3 130.75
R5529 a_2479_9004.n31 a_2479_9004.t0 130.75
R5530 a_2479_9004.t4 a_2479_9004.n0 91.3557
R5531 a_2479_9004.n31 a_2479_9004.t2 91.3557
R5532 a_2479_9004.n49 a_2479_9004.n48 86.5152
R5533 a_2479_9004.n72 a_2479_9004.n5 86.5152
R5534 a_2479_9004.n33 a_2479_9004.n24 30.3012
R5535 a_2479_9004.n71 a_2479_9004.n70 30.3012
R5536 a_2479_9004.n11 a_2479_9004.t8 28.5655
R5537 a_2479_9004.n11 a_2479_9004.t6 28.5655
R5538 a_2479_9004.n10 a_2479_9004.t12 28.5655
R5539 a_2479_9004.n10 a_2479_9004.t10 28.5655
R5540 a_2479_9004.n47 a_2479_9004.n23 24.8476
R5541 a_2479_9004.n55 a_2479_9004.n4 24.8476
R5542 a_2479_9004.n46 a_2479_9004.n30 23.3417
R5543 a_2479_9004.n57 a_2479_9004.n6 23.3417
R5544 a_2479_9004.n50 a_2479_9004.n49 22.0256
R5545 a_2479_9004.n54 a_2479_9004.n5 22.0256
R5546 a_2479_9004.n43 a_2479_9004.n29 21.8358
R5547 a_2479_9004.n59 a_2479_9004.n3 21.8358
R5548 a_2479_9004.n41 a_2479_9004.n28 20.3299
R5549 a_2479_9004.n61 a_2479_9004.n7 20.3299
R5550 a_2479_9004.n39 a_2479_9004.n27 18.824
R5551 a_2479_9004.n63 a_2479_9004.n2 18.824
R5552 a_2479_9004.n20 a_2479_9004.n18 17.4823
R5553 a_2479_9004.n37 a_2479_9004.n26 17.3181
R5554 a_2479_9004.n65 a_2479_9004.n8 17.3181
R5555 a_2479_9004.n48 a_2479_9004.n24 16.3559
R5556 a_2479_9004.n72 a_2479_9004.n71 16.3559
R5557 a_2479_9004.n35 a_2479_9004.n25 15.8123
R5558 a_2479_9004.n67 a_2479_9004.n1 15.8123
R5559 a_2479_9004.n20 a_2479_9004.n19 14.6053
R5560 a_2479_9004.n52 a_2479_9004.n51 14.377
R5561 a_2479_9004.n49 a_2479_9004.n23 12.7256
R5562 a_2479_9004.n55 a_2479_9004.n5 12.7256
R5563 a_2479_9004.n33 a_2479_9004.n25 11.2946
R5564 a_2479_9004.n70 a_2479_9004.n1 11.2946
R5565 a_2479_9004.n21 a_2479_9004.n20 10.4849
R5566 a_2479_9004.n35 a_2479_9004.n26 9.78874
R5567 a_2479_9004.n67 a_2479_9004.n8 9.78874
R5568 a_2479_9004.n23 a_2479_9004.n22 9.3005
R5569 a_2479_9004.n46 a_2479_9004.n45 9.3005
R5570 a_2479_9004.n44 a_2479_9004.n43 9.3005
R5571 a_2479_9004.n42 a_2479_9004.n41 9.3005
R5572 a_2479_9004.n40 a_2479_9004.n39 9.3005
R5573 a_2479_9004.n38 a_2479_9004.n37 9.3005
R5574 a_2479_9004.n36 a_2479_9004.n35 9.3005
R5575 a_2479_9004.n34 a_2479_9004.n33 9.3005
R5576 a_2479_9004.n56 a_2479_9004.n55 9.3005
R5577 a_2479_9004.n58 a_2479_9004.n57 9.3005
R5578 a_2479_9004.n60 a_2479_9004.n59 9.3005
R5579 a_2479_9004.n62 a_2479_9004.n61 9.3005
R5580 a_2479_9004.n64 a_2479_9004.n63 9.3005
R5581 a_2479_9004.n66 a_2479_9004.n65 9.3005
R5582 a_2479_9004.n68 a_2479_9004.n67 9.3005
R5583 a_2479_9004.n70 a_2479_9004.n69 9.3005
R5584 a_2479_9004.n21 a_2479_9004.n17 8.69704
R5585 a_2479_9004.n37 a_2479_9004.n27 8.28285
R5586 a_2479_9004.n65 a_2479_9004.n2 8.28285
R5587 a_2479_9004.n39 a_2479_9004.n28 6.77697
R5588 a_2479_9004.n63 a_2479_9004.n7 6.77697
R5589 a_2479_9004.n52 a_2479_9004.n50 6.19091
R5590 a_2479_9004.n41 a_2479_9004.n29 5.27109
R5591 a_2479_9004.n61 a_2479_9004.n3 5.27109
R5592 a_2479_9004.n43 a_2479_9004.n30 3.76521
R5593 a_2479_9004.n59 a_2479_9004.n6 3.76521
R5594 a_2479_9004.n54 a_2479_9004.n53 3.31388
R5595 a_2479_9004.n48 a_2479_9004.t17 2.48621
R5596 a_2479_9004.n48 a_2479_9004.t1 2.48621
R5597 a_2479_9004.n51 a_2479_9004.t14 2.48621
R5598 a_2479_9004.n51 a_2479_9004.t13 2.48621
R5599 a_2479_9004.n18 a_2479_9004.t16 2.48621
R5600 a_2479_9004.n18 a_2479_9004.t15 2.48621
R5601 a_2479_9004.n19 a_2479_9004.t20 2.48621
R5602 a_2479_9004.n19 a_2479_9004.t19 2.48621
R5603 a_2479_9004.t4 a_2479_9004.n72 2.48621
R5604 a_2479_9004.n72 a_2479_9004.t18 2.48621
R5605 a_2479_9004.n32 a_2479_9004.n24 2.36936
R5606 a_2479_9004.n71 a_2479_9004.n9 2.36936
R5607 a_2479_9004.n53 a_2479_9004.n52 2.30287
R5608 a_2479_9004.n47 a_2479_9004.n46 2.25932
R5609 a_2479_9004.n57 a_2479_9004.n4 2.25932
R5610 a_2479_9004.n53 a_2479_9004.n21 1.07418
R5611 a_2479_9004.n9 a_2479_9004.n0 0.320353
R5612 a_2479_9004.n32 a_2479_9004.n31 0.320353
R5613 a_2479_9004.n50 a_2479_9004.n22 0.196152
R5614 a_2479_9004.n45 a_2479_9004.n22 0.196152
R5615 a_2479_9004.n45 a_2479_9004.n44 0.196152
R5616 a_2479_9004.n44 a_2479_9004.n42 0.196152
R5617 a_2479_9004.n42 a_2479_9004.n40 0.196152
R5618 a_2479_9004.n40 a_2479_9004.n38 0.196152
R5619 a_2479_9004.n38 a_2479_9004.n36 0.196152
R5620 a_2479_9004.n36 a_2479_9004.n34 0.196152
R5621 a_2479_9004.n34 a_2479_9004.n32 0.196152
R5622 a_2479_9004.n56 a_2479_9004.n54 0.196152
R5623 a_2479_9004.n58 a_2479_9004.n56 0.196152
R5624 a_2479_9004.n60 a_2479_9004.n58 0.196152
R5625 a_2479_9004.n62 a_2479_9004.n60 0.196152
R5626 a_2479_9004.n64 a_2479_9004.n62 0.196152
R5627 a_2479_9004.n66 a_2479_9004.n64 0.196152
R5628 a_2479_9004.n68 a_2479_9004.n66 0.196152
R5629 a_2479_9004.n69 a_2479_9004.n68 0.196152
R5630 a_2479_9004.n69 a_2479_9004.n9 0.196152
R5631 a_2479_9004.n15 a_2479_9004.n14 0.0850588
R5632 a_2479_9004.n13 a_2479_9004.n12 0.0427794
R5633 a_2479_9004.n14 a_2479_9004.n13 0.0427794
R5634 a_2479_9004.n16 a_2479_9004.n15 0.0427794
R5635 a_2479_9004.n17 a_2479_9004.n16 0.0427794
R5636 a_3758_2896.n39 a_3758_2896.n4 185
R5637 a_3758_2896.n39 a_3758_2896.n6 185
R5638 a_3758_2896.n39 a_3758_2896.n3 185
R5639 a_3758_2896.n39 a_3758_2896.n7 185
R5640 a_3758_2896.n39 a_3758_2896.n2 185
R5641 a_3758_2896.n39 a_3758_2896.n8 185
R5642 a_3758_2896.n39 a_3758_2896.n1 185
R5643 a_3758_2896.n0 a_3758_2896.t0 130.75
R5644 a_3758_2896.t1 a_3758_2896.n0 91.3557
R5645 a_3758_2896.n39 a_3758_2896.n5 86.5152
R5646 a_3758_2896.n38 a_3758_2896.n37 30.3012
R5647 a_3758_2896.n12 a_3758_2896.n10 29.1073
R5648 a_3758_2896.n20 a_3758_2896.n19 27.9576
R5649 a_3758_2896.n18 a_3758_2896.n17 27.9576
R5650 a_3758_2896.n16 a_3758_2896.n15 27.9576
R5651 a_3758_2896.n14 a_3758_2896.n13 27.9576
R5652 a_3758_2896.n12 a_3758_2896.n11 27.9576
R5653 a_3758_2896.n22 a_3758_2896.n4 24.8476
R5654 a_3758_2896.n24 a_3758_2896.n6 23.3417
R5655 a_3758_2896.n21 a_3758_2896.n5 22.0256
R5656 a_3758_2896.n26 a_3758_2896.n3 21.8358
R5657 a_3758_2896.n28 a_3758_2896.n7 20.3299
R5658 a_3758_2896.n30 a_3758_2896.n2 18.824
R5659 a_3758_2896.n32 a_3758_2896.n8 17.3181
R5660 a_3758_2896.n39 a_3758_2896.n38 16.3559
R5661 a_3758_2896.n34 a_3758_2896.n1 15.8123
R5662 a_3758_2896.n22 a_3758_2896.n5 12.7256
R5663 a_3758_2896.n21 a_3758_2896.n20 12.0517
R5664 a_3758_2896.n37 a_3758_2896.n1 11.2946
R5665 a_3758_2896.n34 a_3758_2896.n8 9.78874
R5666 a_3758_2896.n23 a_3758_2896.n22 9.3005
R5667 a_3758_2896.n25 a_3758_2896.n24 9.3005
R5668 a_3758_2896.n27 a_3758_2896.n26 9.3005
R5669 a_3758_2896.n29 a_3758_2896.n28 9.3005
R5670 a_3758_2896.n31 a_3758_2896.n30 9.3005
R5671 a_3758_2896.n33 a_3758_2896.n32 9.3005
R5672 a_3758_2896.n35 a_3758_2896.n34 9.3005
R5673 a_3758_2896.n37 a_3758_2896.n36 9.3005
R5674 a_3758_2896.n32 a_3758_2896.n2 8.28285
R5675 a_3758_2896.n30 a_3758_2896.n7 6.77697
R5676 a_3758_2896.n19 a_3758_2896.t7 5.8005
R5677 a_3758_2896.n19 a_3758_2896.t9 5.8005
R5678 a_3758_2896.n17 a_3758_2896.t8 5.8005
R5679 a_3758_2896.n17 a_3758_2896.t13 5.8005
R5680 a_3758_2896.n15 a_3758_2896.t4 5.8005
R5681 a_3758_2896.n15 a_3758_2896.t3 5.8005
R5682 a_3758_2896.n13 a_3758_2896.t11 5.8005
R5683 a_3758_2896.n13 a_3758_2896.t10 5.8005
R5684 a_3758_2896.n11 a_3758_2896.t2 5.8005
R5685 a_3758_2896.n11 a_3758_2896.t12 5.8005
R5686 a_3758_2896.n10 a_3758_2896.t5 5.8005
R5687 a_3758_2896.n10 a_3758_2896.t6 5.8005
R5688 a_3758_2896.n28 a_3758_2896.n3 5.27109
R5689 a_3758_2896.n26 a_3758_2896.n6 3.76521
R5690 a_3758_2896.t1 a_3758_2896.n39 2.48621
R5691 a_3758_2896.n39 a_3758_2896.t14 2.48621
R5692 a_3758_2896.n38 a_3758_2896.n9 2.36936
R5693 a_3758_2896.n16 a_3758_2896.n14 2.30199
R5694 a_3758_2896.n24 a_3758_2896.n4 2.25932
R5695 a_3758_2896.n14 a_3758_2896.n12 1.1502
R5696 a_3758_2896.n18 a_3758_2896.n16 1.1502
R5697 a_3758_2896.n20 a_3758_2896.n18 1.1502
R5698 a_3758_2896.n9 a_3758_2896.n0 0.320353
R5699 a_3758_2896.n23 a_3758_2896.n21 0.196152
R5700 a_3758_2896.n25 a_3758_2896.n23 0.196152
R5701 a_3758_2896.n27 a_3758_2896.n25 0.196152
R5702 a_3758_2896.n29 a_3758_2896.n27 0.196152
R5703 a_3758_2896.n31 a_3758_2896.n29 0.196152
R5704 a_3758_2896.n33 a_3758_2896.n31 0.196152
R5705 a_3758_2896.n35 a_3758_2896.n33 0.196152
R5706 a_3758_2896.n36 a_3758_2896.n35 0.196152
R5707 a_3758_2896.n36 a_3758_2896.n9 0.196152
R5708 EN.n0 EN.t0 262.997
R5709 EN.n1 EN.t1 262.007
R5710 EN.n0 EN.t2 262.007
R5711 EN.n1 EN.n0 0.989232
R5712 EN EN.n1 0.365614
R5713 IBIAS.n26 IBIAS.n25 185
R5714 IBIAS.n26 IBIAS.n8 185
R5715 IBIAS.n26 IBIAS.n7 185
R5716 IBIAS.n26 IBIAS.n6 185
R5717 IBIAS.n26 IBIAS.n5 185
R5718 IBIAS.n26 IBIAS.n4 185
R5719 IBIAS.n26 IBIAS.n3 185
R5720 IBIAS.n9 IBIAS.t1 130.75
R5721 IBIAS.n9 IBIAS.t2 91.3557
R5722 IBIAS.n27 IBIAS.n26 86.5152
R5723 IBIAS.n11 IBIAS.n2 30.3012
R5724 IBIAS.n25 IBIAS.n1 24.8476
R5725 IBIAS.n24 IBIAS.n8 23.3417
R5726 IBIAS.n28 IBIAS.n27 22.0256
R5727 IBIAS.n21 IBIAS.n7 21.8358
R5728 IBIAS.n19 IBIAS.n6 20.3299
R5729 IBIAS.n17 IBIAS.n5 18.824
R5730 IBIAS.n15 IBIAS.n4 17.3181
R5731 IBIAS.n26 IBIAS.n2 16.3559
R5732 IBIAS.n13 IBIAS.n3 15.8123
R5733 IBIAS.n27 IBIAS.n1 12.7256
R5734 IBIAS.n11 IBIAS.n3 11.2946
R5735 IBIAS.n13 IBIAS.n4 9.78874
R5736 IBIAS.n1 IBIAS.n0 9.3005
R5737 IBIAS.n24 IBIAS.n23 9.3005
R5738 IBIAS.n22 IBIAS.n21 9.3005
R5739 IBIAS.n20 IBIAS.n19 9.3005
R5740 IBIAS.n18 IBIAS.n17 9.3005
R5741 IBIAS.n16 IBIAS.n15 9.3005
R5742 IBIAS.n14 IBIAS.n13 9.3005
R5743 IBIAS.n12 IBIAS.n11 9.3005
R5744 IBIAS.n15 IBIAS.n5 8.28285
R5745 IBIAS.n17 IBIAS.n6 6.77697
R5746 IBIAS.n19 IBIAS.n7 5.27109
R5747 IBIAS IBIAS.n28 5.23142
R5748 IBIAS.n21 IBIAS.n8 3.76521
R5749 IBIAS.n26 IBIAS.t2 2.48621
R5750 IBIAS.n26 IBIAS.t0 2.48621
R5751 IBIAS.n10 IBIAS.n2 2.36936
R5752 IBIAS.n25 IBIAS.n24 2.25932
R5753 IBIAS.n10 IBIAS.n9 0.320353
R5754 IBIAS.n28 IBIAS.n0 0.196152
R5755 IBIAS.n23 IBIAS.n0 0.196152
R5756 IBIAS.n23 IBIAS.n22 0.196152
R5757 IBIAS.n22 IBIAS.n20 0.196152
R5758 IBIAS.n20 IBIAS.n18 0.196152
R5759 IBIAS.n18 IBIAS.n16 0.196152
R5760 IBIAS.n16 IBIAS.n14 0.196152
R5761 IBIAS.n14 IBIAS.n12 0.196152
R5762 IBIAS.n12 IBIAS.n10 0.196152
C6 IBIAS VSS 2.5517f
C7 EN VSS 3.44783f
C8 VP VSS 5.00274f
C9 VN VSS 5.17776f
C10 VOUT VSS 29.58985f
C11 VDD VSS 14.67527f
C12 a_2479_9004.t3 VSS 1.50187f $ **FLOATING
C13 a_2479_9004.n0 VSS 2.87497f $ **FLOATING
C14 a_2479_9004.n5 VSS 0.01065f $ **FLOATING
C15 a_2479_9004.t18 VSS 0.15099f $ **FLOATING
C16 a_2479_9004.n9 VSS 0.40499f $ **FLOATING
C17 a_2479_9004.t12 VSS 0.02157f $ **FLOATING
C18 a_2479_9004.t10 VSS 0.02157f $ **FLOATING
C19 a_2479_9004.n10 VSS 0.04515f $ **FLOATING
C20 a_2479_9004.t8 VSS 0.02157f $ **FLOATING
C21 a_2479_9004.t6 VSS 0.02157f $ **FLOATING
C22 a_2479_9004.n11 VSS 0.04515f $ **FLOATING
C23 a_2479_9004.t23 VSS 0.09373f $ **FLOATING
C24 a_2479_9004.t7 VSS 0.09373f $ **FLOATING
C25 a_2479_9004.n13 VSS 0.23774f $ **FLOATING
C26 a_2479_9004.t24 VSS 0.09373f $ **FLOATING
C27 a_2479_9004.t5 VSS 0.09373f $ **FLOATING
C28 a_2479_9004.n14 VSS 0.24805f $ **FLOATING
C29 a_2479_9004.t11 VSS 0.09373f $ **FLOATING
C30 a_2479_9004.t21 VSS 0.09373f $ **FLOATING
C31 a_2479_9004.n15 VSS 0.24805f $ **FLOATING
C32 a_2479_9004.n16 VSS 0.23774f $ **FLOATING
C33 a_2479_9004.t9 VSS 0.09373f $ **FLOATING
C34 a_2479_9004.t22 VSS 0.09373f $ **FLOATING
C35 a_2479_9004.n17 VSS 0.94441f $ **FLOATING
C36 a_2479_9004.t16 VSS 0.15099f $ **FLOATING
C37 a_2479_9004.t15 VSS 0.15099f $ **FLOATING
C38 a_2479_9004.n18 VSS 0.83797f $ **FLOATING
C39 a_2479_9004.t20 VSS 0.15099f $ **FLOATING
C40 a_2479_9004.t19 VSS 0.15099f $ **FLOATING
C41 a_2479_9004.n19 VSS 0.6229f $ **FLOATING
C42 a_2479_9004.n20 VSS 3.08737f $ **FLOATING
C43 a_2479_9004.n21 VSS 1.8669f $ **FLOATING
C44 a_2479_9004.n22 VSS 0.02463f $ **FLOATING
C45 a_2479_9004.n23 VSS 0.01693f $ **FLOATING
C46 a_2479_9004.t17 VSS 0.15099f $ **FLOATING
C47 a_2479_9004.n24 VSS 0.02039f $ **FLOATING
C48 a_2479_9004.t2 VSS 0.07974f $ **FLOATING
C49 a_2479_9004.t0 VSS 1.50187f $ **FLOATING
C50 a_2479_9004.n31 VSS 2.87497f $ **FLOATING
C51 a_2479_9004.n32 VSS 0.40499f $ **FLOATING
C52 a_2479_9004.n33 VSS 0.01642f $ **FLOATING
C53 a_2479_9004.n34 VSS 0.02463f $ **FLOATING
C54 a_2479_9004.n36 VSS 0.02463f $ **FLOATING
C55 a_2479_9004.n38 VSS 0.02463f $ **FLOATING
C56 a_2479_9004.n40 VSS 0.02463f $ **FLOATING
C57 a_2479_9004.n42 VSS 0.02463f $ **FLOATING
C58 a_2479_9004.n44 VSS 0.02463f $ **FLOATING
C59 a_2479_9004.n45 VSS 0.02463f $ **FLOATING
C60 a_2479_9004.t1 VSS 0.15099f $ **FLOATING
C61 a_2479_9004.n48 VSS 0.32302f $ **FLOATING
C62 a_2479_9004.n49 VSS 0.01065f $ **FLOATING
C63 a_2479_9004.n50 VSS 0.37922f $ **FLOATING
C64 a_2479_9004.t14 VSS 0.15099f $ **FLOATING
C65 a_2479_9004.t13 VSS 0.15099f $ **FLOATING
C66 a_2479_9004.n51 VSS 0.60795f $ **FLOATING
C67 a_2479_9004.n52 VSS 1.42234f $ **FLOATING
C68 a_2479_9004.n53 VSS 0.3605f $ **FLOATING
C69 a_2479_9004.n54 VSS 0.19419f $ **FLOATING
C70 a_2479_9004.n55 VSS 0.01693f $ **FLOATING
C71 a_2479_9004.n56 VSS 0.02463f $ **FLOATING
C72 a_2479_9004.n58 VSS 0.02463f $ **FLOATING
C73 a_2479_9004.n60 VSS 0.02463f $ **FLOATING
C74 a_2479_9004.n62 VSS 0.02463f $ **FLOATING
C75 a_2479_9004.n64 VSS 0.02463f $ **FLOATING
C76 a_2479_9004.n66 VSS 0.02463f $ **FLOATING
C77 a_2479_9004.n68 VSS 0.02463f $ **FLOATING
C78 a_2479_9004.n69 VSS 0.02463f $ **FLOATING
C79 a_2479_9004.n70 VSS 0.01642f $ **FLOATING
C80 a_2479_9004.n71 VSS 0.02039f $ **FLOATING
C81 a_2479_9004.n72 VSS 0.32302f $ **FLOATING
C82 a_2479_9004.t4 VSS 0.23073f $ **FLOATING
C83 VN.t0 VSS 1.3922f $ **FLOATING
C84 VN.t1 VSS 1.38823f $ **FLOATING
C85 VN.n0 VSS 1.2253f $ **FLOATING
C86 VN.t4 VSS 1.38823f $ **FLOATING
C87 VN.n1 VSS 0.61184f $ **FLOATING
C88 VN.t5 VSS 1.38951f $ **FLOATING
C89 VN.n2 VSS 1.08963f $ **FLOATING
C90 VN.t7 VSS 1.38792f $ **FLOATING
C91 VN.t2 VSS 1.39115f $ **FLOATING
C92 VN.t6 VSS 1.38792f $ **FLOATING
C93 VN.n3 VSS 1.21058f $ **FLOATING
C94 VN.n4 VSS 0.57945f $ **FLOATING
C95 VN.t3 VSS 1.3877f $ **FLOATING
C96 VN.n5 VSS 0.60129f $ **FLOATING
C97 VN.n6 VSS 0.69029f $ **FLOATING
C98 a_2995_7336.t2 VSS 0.11279f $ **FLOATING
C99 a_2995_7336.t3 VSS 0.11279f $ **FLOATING
C100 a_2995_7336.t18 VSS 0.11279f $ **FLOATING
C101 a_2995_7336.n0 VSS 0.32272f $ **FLOATING
C102 a_2995_7336.t6 VSS 0.11279f $ **FLOATING
C103 a_2995_7336.t12 VSS 0.11279f $ **FLOATING
C104 a_2995_7336.n1 VSS 0.32268f $ **FLOATING
C105 a_2995_7336.t19 VSS 0.11279f $ **FLOATING
C106 a_2995_7336.t4 VSS 0.11279f $ **FLOATING
C107 a_2995_7336.n2 VSS 0.32272f $ **FLOATING
C108 a_2995_7336.n3 VSS 1.26812f $ **FLOATING
C109 a_2995_7336.t1 VSS 0.11279f $ **FLOATING
C110 a_2995_7336.t17 VSS 0.11279f $ **FLOATING
C111 a_2995_7336.n4 VSS 0.32268f $ **FLOATING
C112 a_2995_7336.t13 VSS 0.11279f $ **FLOATING
C113 a_2995_7336.t5 VSS 0.11279f $ **FLOATING
C114 a_2995_7336.n5 VSS 0.32272f $ **FLOATING
C115 a_2995_7336.n6 VSS 0.0184f $ **FLOATING
C116 a_2995_7336.n7 VSS 0.01264f $ **FLOATING
C117 a_2995_7336.t16 VSS 0.11279f $ **FLOATING
C118 a_2995_7336.n8 VSS 0.01523f $ **FLOATING
C119 a_2995_7336.t11 VSS 0.05957f $ **FLOATING
C120 a_2995_7336.t9 VSS 1.12173f $ **FLOATING
C121 a_2995_7336.n15 VSS 2.1269f $ **FLOATING
C122 a_2995_7336.n16 VSS 0.30254f $ **FLOATING
C123 a_2995_7336.n17 VSS 0.01227f $ **FLOATING
C124 a_2995_7336.n18 VSS 0.0184f $ **FLOATING
C125 a_2995_7336.n20 VSS 0.0184f $ **FLOATING
C126 a_2995_7336.n22 VSS 0.0184f $ **FLOATING
C127 a_2995_7336.n24 VSS 0.0184f $ **FLOATING
C128 a_2995_7336.n26 VSS 0.0184f $ **FLOATING
C129 a_2995_7336.n28 VSS 0.0184f $ **FLOATING
C130 a_2995_7336.n29 VSS 0.0184f $ **FLOATING
C131 a_2995_7336.t10 VSS 0.11279f $ **FLOATING
C132 a_2995_7336.n32 VSS 0.24131f $ **FLOATING
C133 a_2995_7336.n34 VSS 0.18922f $ **FLOATING
C134 a_2995_7336.t15 VSS 0.11279f $ **FLOATING
C135 a_2995_7336.t7 VSS 0.11279f $ **FLOATING
C136 a_2995_7336.n35 VSS 0.32268f $ **FLOATING
C137 a_2995_7336.t8 VSS 0.11279f $ **FLOATING
C138 a_2995_7336.t14 VSS 0.11279f $ **FLOATING
C139 a_2995_7336.n36 VSS 0.32272f $ **FLOATING
C140 a_2995_7336.n37 VSS 1.58502f $ **FLOATING
C141 a_2995_7336.n38 VSS 1.93909f $ **FLOATING
C142 a_2995_7336.n39 VSS 1.60509f $ **FLOATING
C143 a_2995_7336.n40 VSS 1.26812f $ **FLOATING
C144 a_2995_7336.n41 VSS 0.32268f $ **FLOATING
C145 a_2995_7336.t0 VSS 0.11279f $ **FLOATING
C146 VP.t7 VSS 1.39761f $ **FLOATING
C147 VP.t6 VSS 1.39363f $ **FLOATING
C148 VP.n0 VSS 1.23006f $ **FLOATING
C149 VP.t2 VSS 1.39363f $ **FLOATING
C150 VP.n1 VSS 0.61421f $ **FLOATING
C151 VP.t1 VSS 1.39491f $ **FLOATING
C152 VP.n2 VSS 1.09386f $ **FLOATING
C153 VP.t3 VSS 1.39656f $ **FLOATING
C154 VP.t5 VSS 1.39331f $ **FLOATING
C155 VP.n3 VSS 1.21529f $ **FLOATING
C156 VP.t4 VSS 1.39331f $ **FLOATING
C157 VP.n4 VSS 0.5817f $ **FLOATING
C158 VP.t0 VSS 1.39309f $ **FLOATING
C159 VP.n5 VSS 0.60363f $ **FLOATING
C160 VP.n6 VSS 0.6844f $ **FLOATING
C161 VDD.t46 VSS 0.03731f $ **FLOATING
C162 VDD.t22 VSS 0.01297f $ **FLOATING
C163 VDD.n0 VSS 0.01158f $ **FLOATING
C164 VDD.t45 VSS 0.03445f $ **FLOATING
C165 VDD.n1 VSS 0.20124f $ **FLOATING
C166 VDD.n2 VSS 0.01757f $ **FLOATING
C167 VDD.n3 VSS 0.18626f $ **FLOATING
C168 VDD.n4 VSS 0.01757f $ **FLOATING
C169 VDD.n5 VSS 0.12579f $ **FLOATING
C170 VDD.n6 VSS 0.01757f $ **FLOATING
C171 VDD.n7 VSS 0.12579f $ **FLOATING
C172 VDD.n8 VSS 0.01757f $ **FLOATING
C173 VDD.n9 VSS 0.16525f $ **FLOATING
C174 VDD.n10 VSS 0.05234f $ **FLOATING
C175 VDD.t42 VSS 0.01585f $ **FLOATING
C176 VDD.n11 VSS 0.02496f $ **FLOATING
C177 VDD.n12 VSS 0.0254f $ **FLOATING
C178 VDD.t52 VSS 0.03449f $ **FLOATING
C179 VDD.t60 VSS 0.06762f $ **FLOATING
C180 VDD.t61 VSS 0.03737f $ **FLOATING
C181 VDD.n13 VSS 0.04504f $ **FLOATING
C182 VDD.n14 VSS 0.01652f $ **FLOATING
C183 VDD.n15 VSS 0.02031f $ **FLOATING
C184 VDD.n16 VSS 0.07597f $ **FLOATING
C185 VDD.n17 VSS 0.04084f $ **FLOATING
C186 VDD.t41 VSS 0.06758f $ **FLOATING
C187 VDD.n18 VSS 0.0254f $ **FLOATING
C188 VDD.n19 VSS 0.04084f $ **FLOATING
C189 VDD.t71 VSS 0.0676f $ **FLOATING
C190 VDD.n20 VSS 0.05961f $ **FLOATING
C191 VDD.n21 VSS 0.01947f $ **FLOATING
C192 VDD.n22 VSS 0.02031f $ **FLOATING
C193 VDD.n23 VSS 0.01652f $ **FLOATING
C194 VDD.t72 VSS 0.01585f $ **FLOATING
C195 VDD.n24 VSS 0.01653f $ **FLOATING
C196 VDD.t53 VSS 0.01585f $ **FLOATING
C197 VDD.n25 VSS 0.01653f $ **FLOATING
C198 VDD.n26 VSS 0.10797f $ **FLOATING
C199 VDD.n27 VSS 0.01757f $ **FLOATING
C200 VDD.n28 VSS 0.24229f $ **FLOATING
C201 VDD.n29 VSS 0.05234f $ **FLOATING
C202 VDD.n30 VSS 0.02031f $ **FLOATING
C203 VDD.t40 VSS 0.02945f $ **FLOATING
C204 VDD.n31 VSS 0.07597f $ **FLOATING
C205 VDD.n32 VSS 0.0254f $ **FLOATING
C206 VDD.t73 VSS 0.03449f $ **FLOATING
C207 VDD.n33 VSS 0.01947f $ **FLOATING
C208 VDD.n34 VSS 0.05961f $ **FLOATING
C209 VDD.t54 VSS 0.0676f $ **FLOATING
C210 VDD.n35 VSS 0.02496f $ **FLOATING
C211 VDD.n36 VSS 0.04084f $ **FLOATING
C212 VDD.t56 VSS 0.06758f $ **FLOATING
C213 VDD.n37 VSS 0.0254f $ **FLOATING
C214 VDD.n38 VSS 0.04084f $ **FLOATING
C215 VDD.t38 VSS 0.06762f $ **FLOATING
C216 VDD.n39 VSS 0.04504f $ **FLOATING
C217 VDD.n40 VSS 0.02031f $ **FLOATING
C218 VDD.n41 VSS 0.01652f $ **FLOATING
C219 VDD.t57 VSS 0.01585f $ **FLOATING
C220 VDD.n42 VSS 0.01652f $ **FLOATING
C221 VDD.t55 VSS 0.01585f $ **FLOATING
C222 VDD.n43 VSS 0.01653f $ **FLOATING
C223 VDD.t74 VSS 0.01585f $ **FLOATING
C224 VDD.n44 VSS 0.01653f $ **FLOATING
C225 VDD.n45 VSS 0.08187f $ **FLOATING
C226 VDD.n46 VSS 0.07907f $ **FLOATING
C227 VDD.n52 VSS 0.52419f $ **FLOATING
C228 VDD.n65 VSS 0.01366f $ **FLOATING
C229 VDD.n68 VSS 0.01329f $ **FLOATING
C230 VDD.n71 VSS 0.36378f $ **FLOATING
C231 VDD.n73 VSS 0.01329f $ **FLOATING
C232 VDD.n76 VSS 0.36951f $ **FLOATING
C233 VDD.t8 VSS 0.19478f $ **FLOATING
C234 VDD.n80 VSS 0.37524f $ **FLOATING
C235 VDD.n84 VSS 0.38097f $ **FLOATING
C236 VDD.t15 VSS 0.19478f $ **FLOATING
C237 VDD.n88 VSS 0.3867f $ **FLOATING
C238 VDD.n92 VSS 0.38956f $ **FLOATING
C239 VDD.t2 VSS 0.19478f $ **FLOATING
C240 VDD.t18 VSS 0.19478f $ **FLOATING
C241 VDD.t5 VSS 0.19478f $ **FLOATING
C242 VDD.n99 VSS 0.3867f $ **FLOATING
C243 VDD.t25 VSS 0.19478f $ **FLOATING
C244 VDD.t12 VSS 0.19478f $ **FLOATING
C245 VDD.n106 VSS 0.37524f $ **FLOATING
C246 VDD.t21 VSS 0.19478f $ **FLOATING
C247 VDD.n111 VSS 0.01329f $ **FLOATING
C248 VDD.n112 VSS 0.01329f $ **FLOATING
C249 VDD.t32 VSS 0.19478f $ **FLOATING
C250 VDD.n113 VSS 0.36378f $ **FLOATING
C251 VDD.n114 VSS 0.01329f $ **FLOATING
C252 VDD.n116 VSS 0.52419f $ **FLOATING
C253 VDD.n117 VSS 0.66455f $ **FLOATING
C254 VDD.n136 VSS 0.01366f $ **FLOATING
C255 VDD.n137 VSS 0.01366f $ **FLOATING
C256 VDD.n180 VSS 0.01366f $ **FLOATING
C257 VDD.n181 VSS 0.01366f $ **FLOATING
C258 VDD.n182 VSS 0.01329f $ **FLOATING
C259 VDD.n185 VSS 0.22629f $ **FLOATING
C260 VDD.n191 VSS 0.36951f $ **FLOATING
C261 VDD.n192 VSS 0.22056f $ **FLOATING
C262 VDD.n198 VSS 0.21483f $ **FLOATING
C263 VDD.n204 VSS 0.38097f $ **FLOATING
C264 VDD.n205 VSS 0.2091f $ **FLOATING
C265 VDD.n211 VSS 0.20338f $ **FLOATING
C266 VDD.n217 VSS 0.19765f $ **FLOATING
C267 VDD.n223 VSS 0.19765f $ **FLOATING
C268 VDD.t0 VSS 0.19478f $ **FLOATING
C269 VDD.n229 VSS 0.20338f $ **FLOATING
C270 VDD.n235 VSS 0.2091f $ **FLOATING
C271 VDD.t27 VSS 0.19478f $ **FLOATING
C272 VDD.n241 VSS 0.21483f $ **FLOATING
C273 VDD.n247 VSS 0.22056f $ **FLOATING
C274 VDD.n281 VSS 0.01366f $ **FLOATING
C275 VDD.n282 VSS 0.01329f $ **FLOATING
C276 VDD.t33 VSS 0.19478f $ **FLOATING
C277 VDD.n285 VSS 0.22629f $ **FLOATING
C278 VDD.n288 VSS 0.01329f $ **FLOATING
C279 VDD.n296 VSS 0.01366f $ **FLOATING
C280 VDD.n297 VSS 0.01366f $ **FLOATING
C281 VDD.n299 VSS 0.66455f $ **FLOATING
C282 VDD.n304 VSS 0.08635f $ **FLOATING
C283 VDD.n305 VSS 0.07088f $ **FLOATING
C284 VDD.n306 VSS 0.05234f $ **FLOATING
C285 VDD.t51 VSS 0.01585f $ **FLOATING
C286 VDD.n307 VSS 0.01947f $ **FLOATING
C287 VDD.n308 VSS 0.07597f $ **FLOATING
C288 VDD.n309 VSS 0.04084f $ **FLOATING
C289 VDD.t69 VSS 0.06762f $ **FLOATING
C290 VDD.t70 VSS 0.03737f $ **FLOATING
C291 VDD.n310 VSS 0.01652f $ **FLOATING
C292 VDD.n311 VSS 0.02031f $ **FLOATING
C293 VDD.n312 VSS 0.04504f $ **FLOATING
C294 VDD.n313 VSS 0.0254f $ **FLOATING
C295 VDD.t50 VSS 0.06758f $ **FLOATING
C296 VDD.n314 VSS 0.0254f $ **FLOATING
C297 VDD.t58 VSS 0.03449f $ **FLOATING
C298 VDD.n315 VSS 0.05961f $ **FLOATING
C299 VDD.t75 VSS 0.0676f $ **FLOATING
C300 VDD.n316 VSS 0.04084f $ **FLOATING
C301 VDD.n317 VSS 0.02496f $ **FLOATING
C302 VDD.n318 VSS 0.02031f $ **FLOATING
C303 VDD.n319 VSS 0.01652f $ **FLOATING
C304 VDD.t76 VSS 0.01585f $ **FLOATING
C305 VDD.n320 VSS 0.01653f $ **FLOATING
C306 VDD.t59 VSS 0.01585f $ **FLOATING
C307 VDD.n321 VSS 0.01653f $ **FLOATING
C308 VDD.n322 VSS 0.10814f $ **FLOATING
C309 VDD.n323 VSS 0.01757f $ **FLOATING
C310 VDD.n324 VSS 0.24304f $ **FLOATING
C311 VDD.n325 VSS 0.05234f $ **FLOATING
C312 VDD.n326 VSS 0.02031f $ **FLOATING
C313 VDD.n327 VSS 0.04504f $ **FLOATING
C314 VDD.n328 VSS 0.02496f $ **FLOATING
C315 VDD.t49 VSS 0.02945f $ **FLOATING
C316 VDD.n329 VSS 0.04084f $ **FLOATING
C317 VDD.t43 VSS 0.03449f $ **FLOATING
C318 VDD.t62 VSS 0.0676f $ **FLOATING
C319 VDD.n330 VSS 0.05961f $ **FLOATING
C320 VDD.n331 VSS 0.01947f $ **FLOATING
C321 VDD.n332 VSS 0.0254f $ **FLOATING
C322 VDD.t67 VSS 0.06758f $ **FLOATING
C323 VDD.n333 VSS 0.0254f $ **FLOATING
C324 VDD.t47 VSS 0.06762f $ **FLOATING
C325 VDD.n334 VSS 0.04084f $ **FLOATING
C326 VDD.n335 VSS 0.07597f $ **FLOATING
C327 VDD.n336 VSS 0.02031f $ **FLOATING
C328 VDD.n337 VSS 0.01652f $ **FLOATING
C329 VDD.t68 VSS 0.01585f $ **FLOATING
C330 VDD.n338 VSS 0.01652f $ **FLOATING
C331 VDD.t63 VSS 0.01585f $ **FLOATING
C332 VDD.n339 VSS 0.01653f $ **FLOATING
C333 VDD.t44 VSS 0.01585f $ **FLOATING
C334 VDD.n340 VSS 0.01653f $ **FLOATING
C335 VDD.n341 VSS 0.08187f $ **FLOATING
C336 VDD.n342 VSS 0.09927f $ **FLOATING
C337 VDD.n343 VSS 0.01815f $ **FLOATING
C338 VDD.n344 VSS 0.01757f $ **FLOATING
C339 VDD.n345 VSS 0.32095f $ **FLOATING
C340 VDD.n346 VSS 0.01757f $ **FLOATING
C341 VDD.n347 VSS 0.12579f $ **FLOATING
C342 VDD.n348 VSS 0.01757f $ **FLOATING
C343 VDD.n349 VSS 0.12579f $ **FLOATING
C344 VDD.t66 VSS 0.02938f $ **FLOATING
C345 VDD.n350 VSS 0.01654f $ **FLOATING
C346 VDD.n351 VSS 0.11228f $ **FLOATING
C347 VDD.t64 VSS 0.03445f $ **FLOATING
C348 VDD.n352 VSS 0.07394f $ **FLOATING
C349 VDD.n353 VSS 0.10277f $ **FLOATING
C350 VDD.n354 VSS 0.41351f $ **FLOATING
C351 VDD.n355 VSS 0.26973f $ **FLOATING
C352 VDD.n356 VSS 0.17766f $ **FLOATING
C353 VOUT.t32 VSS 0.03176f $ **FLOATING
C354 VOUT.n10 VSS 0.01519f $ **FLOATING
C355 VOUT.n16 VSS 0.01317f $ **FLOATING
C356 VOUT.n17 VSS 0.02248f $ **FLOATING
C357 VOUT.n20 VSS 0.02268f $ **FLOATING
C358 VOUT.n35 VSS 0.03136f $ **FLOATING
C359 VOUT.t29 VSS 0.03858f $ **FLOATING
C360 VOUT.n45 VSS 0.07315f $ **FLOATING
C361 VOUT.n46 VSS 0.0104f $ **FLOATING
C362 VOUT.n64 VSS 0.03626f $ **FLOATING
C363 VOUT.n65 VSS 0.05437f $ **FLOATING
C364 VOUT.n66 VSS 0.02187f $ **FLOATING
C365 VOUT.t19 VSS 4.93337f $ **FLOATING
C366 VOUT.n67 VSS 0.72309f $ **FLOATING
C367 VOUT.t18 VSS 4.97015f $ **FLOATING
C368 a_2479_7336.t1 VSS 0.01593f $ **FLOATING
C369 a_2479_7336.t14 VSS 2.72377f $ **FLOATING
C370 a_2479_7336.n0 VSS 0.01819f $ **FLOATING
C371 a_2479_7336.n1 VSS 0.0125f $ **FLOATING
C372 a_2479_7336.t11 VSS 0.17038f $ **FLOATING
C373 a_2479_7336.n9 VSS 0.01213f $ **FLOATING
C374 a_2479_7336.t10 VSS 1.10908f $ **FLOATING
C375 a_2479_7336.n10 VSS 2.12308f $ **FLOATING
C376 a_2479_7336.n12 VSS 0.01819f $ **FLOATING
C377 a_2479_7336.n14 VSS 0.01819f $ **FLOATING
C378 a_2479_7336.n16 VSS 0.01819f $ **FLOATING
C379 a_2479_7336.n18 VSS 0.01819f $ **FLOATING
C380 a_2479_7336.n20 VSS 0.01819f $ **FLOATING
C381 a_2479_7336.n22 VSS 0.01819f $ **FLOATING
C382 a_2479_7336.n23 VSS 0.01819f $ **FLOATING
C383 a_2479_7336.n24 VSS 0.29907f $ **FLOATING
C384 a_2479_7336.n25 VSS 0.01506f $ **FLOATING
C385 a_2479_7336.t3 VSS 0.1115f $ **FLOATING
C386 a_2479_7336.n26 VSS 0.23854f $ **FLOATING
C387 a_2479_7336.n28 VSS 0.27998f $ **FLOATING
C388 a_2479_7336.t15 VSS 0.1115f $ **FLOATING
C389 a_2479_7336.t12 VSS 0.1115f $ **FLOATING
C390 a_2479_7336.n29 VSS 0.44893f $ **FLOATING
C391 a_2479_7336.n30 VSS 1.05044f $ **FLOATING
C392 a_2479_7336.n31 VSS 0.01819f $ **FLOATING
C393 a_2479_7336.n32 VSS 0.0125f $ **FLOATING
C394 a_2479_7336.t6 VSS 0.1115f $ **FLOATING
C395 a_2479_7336.n40 VSS 0.01213f $ **FLOATING
C396 a_2479_7336.t9 VSS 0.05889f $ **FLOATING
C397 a_2479_7336.t7 VSS 1.10908f $ **FLOATING
C398 a_2479_7336.n41 VSS 2.12308f $ **FLOATING
C399 a_2479_7336.n43 VSS 0.01819f $ **FLOATING
C400 a_2479_7336.n45 VSS 0.01819f $ **FLOATING
C401 a_2479_7336.n47 VSS 0.01819f $ **FLOATING
C402 a_2479_7336.n49 VSS 0.01819f $ **FLOATING
C403 a_2479_7336.n51 VSS 0.01819f $ **FLOATING
C404 a_2479_7336.n53 VSS 0.01819f $ **FLOATING
C405 a_2479_7336.n54 VSS 0.01819f $ **FLOATING
C406 a_2479_7336.n55 VSS 0.29907f $ **FLOATING
C407 a_2479_7336.n56 VSS 0.01506f $ **FLOATING
C408 a_2479_7336.t8 VSS 0.1115f $ **FLOATING
C409 a_2479_7336.n57 VSS 0.23854f $ **FLOATING
C410 a_2479_7336.n59 VSS 0.1434f $ **FLOATING
C411 a_2479_7336.n60 VSS 0.99841f $ **FLOATING
C412 a_2479_7336.t13 VSS 0.1115f $ **FLOATING
C413 a_2479_7336.t5 VSS 0.1115f $ **FLOATING
C414 a_2479_7336.n61 VSS 0.46002f $ **FLOATING
C415 a_2479_7336.n62 VSS 1.54862f $ **FLOATING
C416 a_2479_7336.t4 VSS 0.1115f $ **FLOATING
C417 a_2479_7336.t2 VSS 0.1115f $ **FLOATING
C418 a_2479_7336.n63 VSS 0.46002f $ **FLOATING
C419 a_2479_7336.n64 VSS 1.39028f $ **FLOATING
C420 a_2479_7336.t17 VSS 0.01593f $ **FLOATING
C421 a_2479_7336.t16 VSS 0.01593f $ **FLOATING
C422 a_2479_7336.n65 VSS 0.03359f $ **FLOATING
C423 a_2479_7336.t31 VSS 0.06931f $ **FLOATING
C424 a_2479_7336.t22 VSS 0.06922f $ **FLOATING
C425 a_2479_7336.n66 VSS 0.12851f $ **FLOATING
C426 a_2479_7336.t24 VSS 0.06922f $ **FLOATING
C427 a_2479_7336.n67 VSS 0.05975f $ **FLOATING
C428 a_2479_7336.n68 VSS 0.15535f $ **FLOATING
C429 a_2479_7336.t27 VSS 0.06922f $ **FLOATING
C430 a_2479_7336.n69 VSS 0.05975f $ **FLOATING
C431 a_2479_7336.t33 VSS 0.06922f $ **FLOATING
C432 a_2479_7336.n70 VSS 0.06847f $ **FLOATING
C433 a_2479_7336.t18 VSS 0.06922f $ **FLOATING
C434 a_2479_7336.n71 VSS 0.06847f $ **FLOATING
C435 a_2479_7336.t29 VSS 0.06922f $ **FLOATING
C436 a_2479_7336.n72 VSS 0.06847f $ **FLOATING
C437 a_2479_7336.t21 VSS 0.06922f $ **FLOATING
C438 a_2479_7336.n73 VSS 0.06847f $ **FLOATING
C439 a_2479_7336.t34 VSS 0.06922f $ **FLOATING
C440 a_2479_7336.n74 VSS 0.11986f $ **FLOATING
C441 a_2479_7336.n75 VSS 2.1749f $ **FLOATING
C442 a_2479_7336.n76 VSS 2.92446f $ **FLOATING
C443 a_2479_7336.t25 VSS 0.06922f $ **FLOATING
C444 a_2479_7336.n77 VSS 0.1166f $ **FLOATING
C445 a_2479_7336.t30 VSS 0.06922f $ **FLOATING
C446 a_2479_7336.n78 VSS 0.06847f $ **FLOATING
C447 a_2479_7336.t20 VSS 0.06922f $ **FLOATING
C448 a_2479_7336.n79 VSS 0.06847f $ **FLOATING
C449 a_2479_7336.t23 VSS 0.06922f $ **FLOATING
C450 a_2479_7336.n80 VSS 0.06847f $ **FLOATING
C451 a_2479_7336.t26 VSS 0.06922f $ **FLOATING
C452 a_2479_7336.n81 VSS 0.06847f $ **FLOATING
C453 a_2479_7336.t32 VSS 0.06922f $ **FLOATING
C454 a_2479_7336.n82 VSS 0.05975f $ **FLOATING
C455 a_2479_7336.t19 VSS 0.06931f $ **FLOATING
C456 a_2479_7336.t28 VSS 0.06922f $ **FLOATING
C457 a_2479_7336.n83 VSS 0.12851f $ **FLOATING
C458 a_2479_7336.t35 VSS 0.06922f $ **FLOATING
C459 a_2479_7336.n84 VSS 0.05975f $ **FLOATING
C460 a_2479_7336.n85 VSS 0.15535f $ **FLOATING
C461 a_2479_7336.n86 VSS 0.03359f $ **FLOATING
C462 a_2479_7336.t0 VSS 0.01593f $ **FLOATING
.ends
